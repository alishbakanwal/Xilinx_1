`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxZhNmo1lcKpLYPA4vXVI
shhj9wquP/jqwNK2XQFYkOoko3u7cVusEV500SZDkSc5oW7XJ6xG7dtlrQuh5jyV
NaKryVeFowXf2LTRteboQ1HsrCRICdpR+qyU9JBg8lRS7LhaqJq0r1EeFJ6W8xof
io9ggEvdWvPGGpZu0hv/fykuRWevDCC5ITcx2GeHeHEKpEsqqBGMUOEyv+MRRdzp
pakAIldB2MRGf2CJqC2Lptcdxry0PQDQHmCsrQi7VxDGdPQp9iq+e6r+wXSqJb7r
yzFcHXII4N4IlaZsBomALCVnsBxLyx1ilKWXsdwOSH0IH1EjTLIqxSx2pJBfkFRr
xQIDAQAB

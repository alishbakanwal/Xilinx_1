XlxV16EB    fa00    15d0F��@�Z&j�Hn�'���?x%0RC������������ �`��U	���Ș�I�F�)Y�g3�4yn��5�/��%���`;�g�dp���2!<#U������\����;��4�E6o��X�>�(�OR�O��
���-P|(l�
�#H�$����(���󐶃|����lg$a;��X��*��&G��R6�Jqz�����n+������td��6OS��Ֆ���/�z��2�����t��o�K�Y�k1�.�o���/?�Ҩ"���7�������<� |P����e\�[�'��i�*�����g܇_�]4���"�~�7[7�K��6r��x�Z��ϓV,c�ÅeɆ��p�d.��~&��8�w<1YI�l@�d�n�nɾ����u�{�$/�E='�_�̹;�Õ~�L��9�n:$�oX�#̮ͤ8�́���*�Dm�9� z,�͠@Ε��p7<nY� ��_5�.��A�h�|�q�z������4E;�b7���(�Zrԓ���j��T�鳨� &^3 [���Ub-��XTs +���z5��7��NM���\�}�x۸x��i��/7���u�"Ŝ�B���'�f��6�#��2��m�%�h�׶��G��͈��5��K4�!�c���E�`��(�G�FM2m�Hv��B���x@p� �z��&'��Du���=}.�8����O�ёHP��,�����
�gA�x���J|Jc�ۋ��E�L�8
r�=0����`>
;t��\�bZiq����@(*����G�_�˕����/J�b58o�=s����p�S��(z�;l�
>�i��O���F�(f��S=���U�F�En(BQ��}v/^�ǆ���	V��\�C���=��F-�m��*iy�:~T#
Y!�9��-Y��@C܄$����ʎ��Q���}�
��li�������F-��l��>[��iu�D���Hd��7�p��w�k�
�S6�'c×��L
 ��s�}I�ƛ?�?���O,�nõ���ʻ �=���y�*�HZ�W��oZcù�@�
�π�"W�09��E����X���ǚ}#���WB�E�U���x��
��q-y��%N'��m�qk|w��7hz�񀍡��e��Z
a�Ǩ#:�S��Z����؊���:G�A����s�:�?����D�S�Џ��K�M�zMv�8I�H\����DQu	��
M�����7�u�(ݺ��+��R_���g�Y��
���`q���ʶ|���]�p��?YָȒ�}���l��&c]��B�v$H0�ܬ��zl��h�ɗ�٦�<J�	]Is�]su������8L�~!�&��ndpU�3�˯ȑ�a��A���4�K�8��`'M0$E�����\o�[���l���"�ts��r�:#@A<79k_�[��'�_rH��7˼��x<}�L#>Ǡ䂶���ݎ�P�	�q�8��-�7"0k���Cج�Ǩ+�{�x����mSC��Eo��a�}�q�b��'l6�A1�dD�M�GN��g��CP>���(~BH�VBCd	���Clv�5?��ܳ�}X�z3T�]�i8o(�yS�S�!Y����ٵ���L���ư݇A���Ė��9���kwe´�bu���b�n�̀��u�܆,�X�QU�)��t=T��L`KjѸ�a�ۃ7��PS-��_�������+�:W��q�ea󊳥?��i�%�w��#tt҉8te�~"�p�����s^�LmӲ�,��0�%�H�A��P���{��uՍ!�q��4����߆��e�aYՕ���4���9�~'�xp3�+/1A!'Y�fH�w�Esy���5e�(�4�� �?x��#D/��[ƃ=��B`�T3r����ny�}��x��N�!WzC�x���HC�RRξ����}nGh�,��o����6E9=n����,V�e[*��[�	˷,����Ve~�x������8��^��C"QY�\��5��@l9��!13�]-r���hEX�$̽��׸тb���{�R�c��<3M�5�i�� ���[�ؘ�v�H�2:��N����O���!׉���9(nC~^�Z��/ ��c3j�M�3HLl[.<��'e��F�j�^���c��8?��{�'�;�g���ra,�r�����^���������C���fY6�	�
����yϙ�����O�n����ќ_�d[�;�JJ)ǥG�<�("`�o�xc�}�u�ǔNՎI��")�d֪y�f� q��A�P
9�~R�,�+�	�����WELtF���[ ����~/:3-����iK�<�)�:�?/�Gw�*�&o��o��/�T|	Π=�\8�Jq3�g�l�&}<@b	M���+)�d��"���$�5?&�����e��~Oդ���=�!xS,I��V�ʱ�06�?<�3���X����4���Z9��%���t�*�2�d13&��^>��mr�jB�w��J���S��}�];[O�Ԭ�c?MXub�;#r���,����U�����^��B<���V���A��[�O�P���b��ǜ���ϡ~\]C88G�KܯeF���-w��CՕ-�٨yǊ�������Ux/B@x���ᖻ�<'�G"`*�?X�p��J��X@q�i!;;i�៟�1�)�E p��kh�����a�AnL��$;?��٨4ρ`��;����W}ͥx��t(Y>g��ޅ^Q�7�hh�����$��!�0�t�񪋡��s����U"^�����H9:#D~X.�U�x�K���>�m��\r��h�]5�?R�Ե4�Ȟ~�R�e�Q���r��]Z^����y��w (�tio#��P�v���v��#aJ�w�:P�?q�0���;Fn�I����fv�S���G��-l��q7]G!���� !y���ç�]�]�	{v����X�-���?7��<����(=L�]~*j�j,�C&���J״*�=>S0�D�{Ak����.��z��45�`||��k4��8��2�A����U�݈��glvJ��"���:�0��AvfR�)bs��p�h�Ԫ�Y�(���!�#sf����xaWE�X�	P��ۘ���ʵ�Icd�3����{}r�y� �嗥y�D��z�VZ�L�?5"��?:P�(�P؈�1J(-i�P�B����	o��E�q����Ӥ�_�l�6��#��E���`T����
գ���Z��j�Ik=Jӎ��X�n�wx�:��K#�:vo@?6�&-C��e�d�8�5*DDc�?�o�\� �����߂*�p��?sb�����%�O������v#1�CTG��L�~ב�|s��:cUt
�* J�cK��d�N�}�E�8#��9fI��Y��x% �s�Ւ���{�𓻳T�$, ���V��w3���Ѳ�E����	?ݚF�ϻ��I��2#�֯��o˴�t�}7)�����^=(���Qx�'1�x���Vǩ8�ijW��[I�<�?��&\-��W
J��m�ǧ����
] T����10����%�§�6]�w.lY�0��֏eL���w��V)�3�B,U�G�V��:� �������ď�ӻ���z��C��x�4�T,�-s�Y�Pd�61�����SUhM+\*pH(m��r譶�"����������>�9�t�L�dz|���s�a���2?��m|´�����}�~O�L΋�L�����"�;�m��I}�P0�A�2-ˁ���Pq �
��8��Nꗴ�o6�a����ր[�J���-�f���b�`���n{�V?.��y���Ջ:�ӎ�D�qu�Z�lH�-Ck�t���Wl�!��-|+����E��ˇ&�~󋝀��T��Uy��_P���"'���lTU��ùS�ڧ9�XP!���_��;��xM�z3ZD�M� ��`�`��k�2k�`Ԅi��s�+�:IF��9_W�w�@c���WJ��/����o&P�"�M�NǓ�؉�gW�`�9�uAm�����Bd
'8�
��kL� [��_�K�۸��m8D�|�3�.5{�9q}��	:v�[�n&!}w��W!���A?p.�j�b[7�$U����r���E4�zX��P9^�la��4���%Js��2]^��U~C.�U��On�����\D�{�K6q�q��(i�E���]ZYj٣il�+������v P���9aq�Z�b��2�b��������y�=���YG�#U3��[���l >ұ�d�h�o%��W���2"�**�
R@�Q�Սt��j����lrW�L�5�5�F;��E���Y���i�IAN����F��M��dx0���{� ���|8s�����&��� aVSg�D!ȸ<�1��S��-���<�kb<Hd�P�.�7�a�A+'a��;�����ԑ��VY�#��`��c�������4�iKv�
����&��UY���9𲲾!2)-�˒��:��,n��<=��Y�RvN�$[�O�d4��s'�s�׾F$4�)"���J����3���vI[ ���.���G�q/��PS�!��0](�۝[�D�y%�+�8����9k䩶�X�.��uA�R��{C����i��(�����2��ɠ��Jݸ���%n��z��qbL�~�*8�X�xun�#�|�x���f6ٮ^ݔ�;���V�^L{\�x�AH�O3��v��Z�VՂ{[�ל�nZĝIE�:�������oV�_�����4X���1��I- _��=�=E�!��ᷴ-mB�(~�5�M-�M$d����[�Y^/n0�(RѵFm6�=^�\�����QB��r����C+q��2�蓾���A	>�>��I"���or$��+��D�1���#N^T_aމ��Q�{�C}�2���t��L�@��A���1�ōC{ݨ+=����b�ki@�&g��fk������0�n���c��g�KWn��2"�B��K��-�:�\f|�~���hC�+~p�z2�V�2S?ƨ�yx˚^��׬2z���)��}�՛�W5�(����CFP:Q��b����t�y�N��L�����ؔ��i��@��J�ol�]�U�)���Ȋ�w>C��R'�iQ��K���0�,���jLy�C�Z��A��`���"�oY����g�oy&��:8����Xb�7�g�+�؇Kto��RzR�~l�{��v?�撨+>b�썚�^�h�Dr&��B��q�Zy��2��é�� �<��2OtR�|�gy��4�
Cϟ�)v˕+�+9ʀy�~��젍ҥ���~B��E���G�^���{���+�F���x3�&�Y�H�S��W�7���L�3~g���>��BwxǄ}�_wc�9�~3�ڵѼl�
*�_�U�E�C����'��CV�����.��xY��U>�P�-�Wz��SC~�_�$?Py�)vy���L����zwV��	����/d�hY]4ӥXlxV16EB    fa00    1500fN2@�$
vb>�l����oi�3�� �򰫆�C�m-Q2��<&��a�ů����yp����Ue�Sb�TEӽE.aBT0��h���L�2�s˽U�����4#.�����?��_'m״p��NTww]l�7S����$��$���l�{�J-�}��2�pi�y<����~��v��QFS�YO�t����]i�5Wm6��V�@�$�t�:��F;"K�Y,,��7�Mu]�]�T�PQ\=��+"#�S�Yꀯ[����������{o���x��Ko�g��3?���k��磪g��?�[E���duG����m#�ц��%��l:.��?Vg\��j�XDcn૙�Ef��࡚ȍ��!�`s�0��l̦�d�]�7�!�]-�i�njm��#c��D/�O�1�*��f�1�$Ԅ��g��7��[Zx��9�����"?��O��,p�ELr
=�U�
�5�=2��Q�M�G�Μ�A�f5�T��
��Vt�:��!�zT(�8z�&Zq������K��w�.������b]�\��������V�f�(d���0Z�MfQX�)t6�^ҜJ��c��z�M�P��;9Q@/����ˎ)9 �Q��&e��k�-Ri	��!��Jw����*S�8�q�B�6.P��S>�|��h����4�+8��`��!�	���zW��.Q��;Ƚd�肝��}�C�q�7��3�छ��ɦd���X���΂��S�LM��߱�������8��dUY\7��
��'Y��{+�)�s�q,oDe��;�J�Wƿ��I�^����������Y�bD!���,�r��g��dBx�>6��[�Nbj���ZG���Y8A��7~��I"����������q� ��H+�{�c��0ڧ�p�&c��c�8w-��g]Zb©�&j�z옶���yp��a|��>c���@xl��b�M�^��p���ؕ�1���ς���\�Qh�67�~��B���f�5�=g�0�5�դU����?��g*u��f���f�D����o0R�څ�?uy]��5�8�G��yвg��B�����{�V�3ո�̋k��F���O<�b��g
^�#w�5{���m�i���J��N+?;1�F�T+I������=n+� ��^�K�x_�}X���
i���1������C^�)�M6 �tS�L*
0u��luR���N��^�z(X���<S+ �
�G���ٻ�8:��pK��<��h&N���
9-�@y�n�f�D��H�V�w��/Ȫ��[�'����i��Da�+��c�B���V+i�d�-qUC�(I�~HԻ��%�^R�oQ�E*�{˷���<cPZ��^�(El��13c���nV��Fy�LaLΑ)���++kTsG+����)}��C-i����7�*�.Z�n:�C���w-߃�I�ϙ�z�������\	����%��6�N���ņ��s��X `OQ5 �����8�sa�\몝>���o[-/�2���W��� ZpB?�]'���/����5�bbD�)D,V{z�y�3�++�θ�q�����sq9�~�D���	u�1��Z�Lo���o� �x���&����X=.L�
�S�}���a�����r��؆�|��$k�:A6�\6 X�b�[#�4(�x�MF5*6����v�x5�	��
������c˖���%�TF3M�w�bO��4d�^񕔼p�Q�M
�9����H�h]���c�5�YCV��:�Ȭa����V&D�~)2�����<�)�+� ٷ���4��Le�� sH��^e���ȋ^���Qx@�F��ڔ���;��������x���0Ra�Bv�}f85�cx�&Pe���E6P�	E�Y�׻�8�Z�s��V��_��W7��U$(Q����SdY���{|
Vݛw�w�(X�P�I������W��������T�؊'��zK�������#�p�d�謟�_"����W���܋Mux�2g�7'ip]�g�_��bo��ٔJ[3�,�,��6�e-ϐw���D_/�̡���J�����=/��گ��b��YN+=�#��o�d�>���у�<�9/.s7�FyQ�~���;\��\�S�5����,�-����L!��)n{��<�{yL��+��7~E���vc9�".K|�l�50��z�W�u��P���7��v�ԍW���Q���P�\Y�U��*��R��B�̫���_��8��ei���`�ث��i�͎�W�=@�:���2����p��iq�;C���.{�g�=kЋl���k�	0�g�"V/w��������*M��)�@T�!a>rF�����yHHSإ��aToZ� y�͍��섒a�4 "
:����1�V8������q�6��	�3��������);}\9W¿s��J(_�
��E�L�p�����QäY[+d�,?��}H���D�FrðD�$��<��c�B��Z�ӊ��>�b�>Y���قG�T��	�>��@Yb�IJ���wT�1�?F����ɀRB;��'�~�䎊��<[�-�n� Ll�����,����9n"k���U���d�R�cW��m�
�1�<���>�Ƀ ���Z��9l�tˏ�������=�v�M��@�����5�K
�uF@>�K���qF��q��� �K%E�!�5���
&(�>{��� �:5n�H��gE^0a87O��8�%01yo<o����	O���9ܨQ���/b�u�?Q$LО���ޖ��pƯ*������a�^�0HpOϊ��&���[^Y}���+C�%R��v���^��S<�B��+�t��r�K&�-\I�����s����� 0nШO�D*@���4Р�����eſ[TE)�G�qǥZ�����1������&e�(ϥ�
�:b�2���N?ĐSj��r6hnYs��lc�RH�Ou;�"�g����Hv�� nN j�7$�{"�U\�۪��ʏ��a�����}`g���C ʊN��֊�׿.+*���
��,�l�s��xNƿ-ȗ5u[�e�g0P+*X�g���nܥ�ݪo�(��"�+�����F���BϽ�K6��اg8>��*|��Ĥ,0����DT�n��Q���Kl��ϸ,�ab�)��\/nb�
�1��_7�[]N��8y�.��	�&��4���K��l��E���Ñ�S͏w#��U�;;�c��9E��F��څ𿕟{,ᗤ�t�\�؅��)逸�x�؛#K��9!	�n�R�f��7i/��#��}����`'���5��x�Q�V7��V6��Dԙ1�U�%���k����D�ؘ�}����Fl��LG���`�ܕ�˰�(<Nچ���d��� ���IY�˯g7p�e3^W�¥�3�Aj���?�2	|�Q�Cάf`Q9D�L��qc�:�K����M?����x5��+�[�(����AT��o+����c�i��{��I ���=a��������]j�jm� ��e��M%���&3Y��Q�(��l�z.W(�-9p�0�m)�q�'�ə�Յ����H��RrU�;	�����������,�_8�|JH�_�hǼ�!���a�U'�4� :*&'A�]i���3b�T�a��s�8x������U�>]�'���ΘBo���n:�3���s<�AGL���v����Vݩ���AV��lȜ��!0ʶ�P[] �k���ly��2v�
9.�u+�qư~�`0#k��O�Ӊ��A&��-��$�g7�҂vڍb�s^�y�`~e�l��A]��?���� g较�z�G�e�Y[�pȩ�	x� yܝ�7�ᰌS)����x�3��	�a/�^RrL�>���WQ����-�̈�m�cc�����J��Hn�
��=�F�ժ���ά��3�{߮����خ[n������,F�g�
6����en�x"+Zq7�y��|X��b�:J�{��]�X�S�#�sgN�x�љ���Lh�!�Z���/q�-H��k�s�y��|K�B�U��p�ʠ^��9�^��h��3��]
��]�������	:^��^_�-cu ���2���H
���T�U�i�!gmO���tUڒIKc� �/�p�
���%��>�j��&�B��e[�l�jk���h~#��.H�/����$�jE�N&J��	'�^Q;�_���9	�52�]�_���~>w`I��a��$�j^��_47��K
�"��Uց�FȰ��h'��M8O�� ��=Z��"\o������B�h�VS�+UE�p� �ON��Ԍ�� 6e����{��0*�)_W[���>�Է�ˈv��po�����e͘��'��Q�	@��]�5J���}�M(h�^�v?e'/�������ϔ���"q��t|�	���ɜ�f�v����0��P�#1D]�S�A�܆If�w��j���h�~�,#��<�d����^܀����#,W;�S�%s�8��/BQ$&������,2'E0�8$���B㮳!L� ,��"���~���fyc@X�8}Y@��CrhWG]=i[/���Q�8%��O��zCЇ!�D�*���|��L�A�}&�A=,~�+�U�MRn*4؀�������5��2y2&[}Q�A��o�d���0�J����"��i!�u��ꖗ����k8����[��H/��I�m���c�����qB�T����9�Ss/����O���m~=ʋ��{I�>�r3�[�$Ye�)�T��A� D��EK-1T=����ā��wH���\��۬�:�T42����Q�����5mtP3���D�����H�0���&�V��31vE��a>���Z����������갽�������J��EP��q�MP�xbk������P!eӲ�W���skW�{��y���[^	��pm�D�4Mu��6c��_${
;����C`U�o'�"�[~�U�)/�Y�,��!��`�˺��&a�@[?�
fJJ���Qd�~����1mF(L�{�Wn��W��|n<���"���H��w�D�·,��LB^Rz���Q��MH���kLa���$��m�
����iY�0�&Bv��R$��zN7P���P�*}�-EW�m$���i	�a��,S}h�c�,>��.�(H�����v� �@L8�F@�)��n��5��v���6�ӕl�Y�������b�7+]��$��׉V=�����8ȏ��NW%��B�km���f�,T`􌳼�&uNXXlxV16EB    fa00    21d0߸Q1��oGm�y�'�^^��:/�f�c6��f���2��L�ɍ{��s�=��
��GEA���ٙ��)���`w�	�p�s0`Q7���u˻������dV�~:>T�1�EX�a�l-�����;j���N���j�5����4ƠB𕁢���%�/8�R��;���!��o�գ����fp'_snK�aAӆ�Z�v�-[s���h3�gS����i���R���
_'ߡ�$���^tF����p<�ȐM�u*�P=l���/8jj��g��s.����q���J
�ǹv:n�W���Hf4��(RE�w�mEhցA,v0��ɏ�8j��7��!*���%HVJ Iꑌ��I��*�	{ �o)���Z�w�R�v�KJ<�{�tk��K�����i�Q�����J_ �e�.O��p/9��΂��j�C�_�e�/��|N�'�IhiTj�� ?-'���)ߒf�{����Lq���+��a΂�cr5���Mg�}*|q��CE�~���E���|1q9:�F�~�>cN��	��a��Њ�uL�RS+��fW�.�Dmh�
����2s4k�i�;e!|;���T��"��،����"�R�<:A��e~�����F�0�N.���v��DZ�Q��p+����{�i���?�l<�.�T�KW{���#=յ�J�������C��9�u@b>�sy���o9�J^z��$�re�0v3�65���ц�;1Hdp��F�g��BP���M�;��"麖_'/]$�	�<�Ծ�w��BMֵR�q�ǥ�Po񣒑N�>��ڔ��92��L���Z��ГY��ܦ��<S�T���G��@ܥ"�ǝ��{(9��ܥ��6	���Q�jJ9좬�&bzT�	�ĝ��S���A*�]�U@��7�{���j�"L[Ϩ��x��#� A��d��P�2�t 
}*ٍ�S��NN(cE;�;�3\�Y>�e$i>.���M��O�玁��w;P[&�뤓�?��f�cZ���I��툅fPL��!09b:�:���q|�i���9	d�f��QT�_6���wԓ蔧*����\��G/�R��_xB\��;^����y�Y(9�����{��`���Ʀ��	͢�����1տ�1F�n~�M�������cs��똨�+�9�yT����V�^|�X�S0N7�pݱ�3�̕�Ȁ�YZ~�B�|8~<�}_���L{��6�����|�ܲ��F�M�4�фRU��c���o�>�-�O���0���
|�_PX6�&ɕ�1�"���e�3R����|�r���/��$T��[�~Rw�(��}�]?z�5F�t��S�h�a<�&�d�6�3yj�X��5����P_%m����F\.�M�ʗ��Ӛ�t06u�QI�B!��k��2��{1��0�̊ hp�V�����'+[8 �FK�][|�r��UBI�"�9��w ��ӫ�E��BR�ē2��R鸺���*摑54�+�6���ч��dR���Ϸ/��zR���	��bK�N���M�OO��g6�y��~�b���]����@+����<��8�><��
�Xb��و�g�R��ϗTq2��C���)��pW%4k��j'�h70��4���S"��iH��k�<��1��nk�v����ب�C �|h5}�HI�)c�߮�$��*��4�~A9�{��N����S�u��F����-L-��m���cEpN�72ݰx�R$Z���1K�4޻�	b�S؁ d����|���IA� �~O��果EL���-�%���ڛ!h9�=�b/ǩso�g�6>}0��������6l�LVZZ U�<���G0��.�b����v�9��$;� �e� �� �s��/��| S��ze"��HuI�nʼ���*�p�}����R�^�q���y��v�X�Y.���$mP&s��sp\!b��l\}?֪4�#4y���	��N#�т�91QX|�L07x�����J:uw�ؾ�L��#IJ`P����R�_�"�c�+T��0;,��+���݁�8����#�Q6H��1�5v|d|-�"��S�6�{^P�Y='���X�D���ME6�g�����ќFH����T�%��-ۛm�����X"�,-[�ֻ�h%��-��	���/zw��c��㟍�n�X=�u�))ZZ���_=�vI�曲�9���WI 
��K��wPI����/�����7��f$;�*2f�eUGdvQ�e�p(*��ֆ)�_Q l���jķԸp$��#C��~���S�mÔ��b�A�L	�1w�V�t3�ᆬ�n(�h���ޜ6��2�W�Ӟd��X%{���ߴ�(���$,2W�j����P�,H8��Am}�i�w3jb�_�uMD>��-��m�. ��+֝�ۘ�<Hu����h�e~~�[2���LD � ����uCN�hJ�e"�Յ.e��3���rGߘA�y���7����W�▾�`:n�9���Gt%쇢=1���� Jhڨ�yN�9�3<6#�o�7��8���8C�"aZ�+ ������O��$d(R/.��F3��Ui{�x��#T�09�Y�K����N�0B�sX�hx��U�^G�:Th��'83�#P�0W��� 6��jw�Vp2i�e]�Vzv[� ��:�(�<F{�
�b�e�=	��H��h�A��jF�hGU�����V3�r��_���������
C>����3U�I�j�=����'t}��T��V7����;;�( ����$f�d
]��؛��7V�7E��r*�-��X�Q��%X�m�K�;�T�kJ<��I�;� ����U%т�R^T�r�y��[��x.���y�kC�+��-𜺄)+�&��}��������>֊�n%���$^��W<�߶c�Nb�B�$+����ΐ�>�j:[��d�]J_���OT���p����
{=���L�ĩ��څ_Z��ʂ���B�%��&�e�n7W��e��^]I�E��7��ID؈�,hM��pw������hNl��<8�7>�m.{��F/r��RZxy�'U����Ha�`Y��}�����Q�3�&!%� �5:����as�A}%fa�	����������F�������I|�������T�6�OוXr1����
�2G��(�p"ol�^��Ԁ$G��Г�Y鷈��=�)��>��Q<�kŤ�!)�N����f�gA��7|�Rڧ���G���$s�:�g�͝"�r�gB���0�Y0!�s��΅�L�׶gd˩]�W��7د�bR��$�1��3�@6��r]5FFo���O5H���J�=���&`rv��I C`�XQ�xK'Uy)5 9y�p{��D�b�^�v�=`�[\�
��1@�<��N�7@���M@g��OC��v��_�:�(|����,��o�2cR�c�7ݟ���@��ʗ�B8���v���o�.�i��k�����på�~�t)ˮ�����b�xsjR�צ����2@ࢨ�hTG�J�T���2��ͻ�?�e\ؖ8��nI�v��`4���_@]^)1�XI��8�L�_� �q�}��y�<҂
�ޏ���oU�+��>�^���1̏����{Z
 �5�vNXi�J�}I���?���,���[����T-�)��E��N�V��+�ǒ�����Y�8.�'�1q�Ӎ�E�n�
�6���=����f���V1B)�Zoj�+O����<W�$��=��$e�Q˻'?[�G	� ��T�(���[T~}��W��߈R�e4	6H���Vg����4��&�_N"�O��Z���`s�GՐ������>:��/��aX��s��0�/S-0'17U�L�V�[01�;ui�5����ZҶ�g���h�X����ٺ���0Ky�P�~��J��=g*���Y�:�6��ͳ��V)l�d���L�-g�`�Ŵp ��pFF��'Ŵx*����A7C�<�C��Ӝ�Iw��TX�٧��)'j��}��P _��w
vΩr�u�+�O���뺫/�=��L�НFp��+�q��}��F9L�.��D�.muN��g��3���*���nu���n��L��kw�����;�Z��Kt8���A�}�kbf���s�n��
��,4CF]m?fq/���1\js�,����Ld���"z��<��܅�����\��X�ICn'��-ՓA��g�FO�Z��K�E�q���9��NІ�>+�M�.r>]?s��lb2���o�-ѧ��l;}�~�������	�������_LB~�Ȧ+��?���'/P�y_��<^��_�۶Rx|n�H?�Lq�붤�3B֥	��.�a�˙�����'�Z�ɡ� 9�`h�s����qK�u�a+��Ph	��fTEM�����`�b��ϗA~Rw�w,���J��8����[�'��p��H7Iz8<"ѵ#D�W�Z���`�kH����(K(d~� Ԗ;�}ڒ0��̪Bn�u|}�9�2�-)
=�w�Ȯ���W�8&��in�3�
v(�TE5Z[T	���j`*c ��3�7�S��N
�>��A�����+�4��1��{�k�|y�)	�%�u^�g3��B�h�Ø��Ue�`�#�L� @�!�g����͓T#b�paH�v��[�Ys��n�YER�t��L���<_ԏ���7����ވ�zwar�ϼ��u�ZÓ���T�/T�|!
7��xA�@o��Ҟ�v�D��ly�"��IW�.�ֹ���F�vdQnse�X0ᵣ.��u�����@. f�D�����]��Қ�?� �>y�{�� �e1Z��w܁�`C�y-6.���J0C����/�b���h�M�&�W
]�Y��]�%�tǪ����<0���AvlߣF��0��ͩ0������|�^m�es���eX3|��%�ח[��<.Ł�]<�X�ڎ��I;�y�|�������]+#��L7@�z��H����mV��"��N�v��]�^՝G��C��;���/�OJ�3��@���������lt|�]��t?�N5�"�.\�����Vn�4f���u�"0��iw�t�AH�5d�����Xr���i�s�0.?3r�����vT��[R�h�1^Է����T"��W,�;9ƍ�9|R�1��L�_�m�y��K1����{��Ĺ2	czdv������c���#=w���+,�D�y�i��a���Nl���t�tU��#���!�Ofa���GuQJ!���&+b��t��QƂ�����\�zF�I}�B���k]'ajҌ�|��V~���@���%"���2%Ƹ+�x�������zcfƤ��X�]3���8h����a�_,��W��i߁U�=�3_
�gTŢe�.&:P֢n�Gf?��ܱ����ɵC�i#Z�%WV����i��<�=J(˅���q),_r���z]k	U.ϝv���+C�/��96
�UZ�牀݆����UV����w	r����M*�i5��\�q�jr�`ŽE߈���6���#
+���-1lq�ԙ�SS��uT�
����� ����P��j��j��U���'�a�V}MO�E;��=S�|�U��UL�c����o Cޕ�1�y��r���������j@���~<G})2�G�ȴ1u����K��|ⱺ_e�$�?���h��J@�xC����!�ȋq�(
����m�ـʛ��<��D6_�T�z���>��T���Zf�L����gt�ң`3�}���<]��}_��	$퍘�#zz^_�ލy�wa��sUlJ��E3��3���aa����2{B"��ޔ��cn(GD~쟻�0j��M@�[�N��˜���H�rv�Ny��7[������!�U��o�����Ӗ0�OWMq���CT�)_ݳ�5l����u��I��Aq�	�6F�o��e�έ��P)��.F��S��G�Ss��pA	I�d�E�8ĲA���Y8�.�Ӊ`C&\9�+,��l5�I�/ ��+6�)�G7�b{�YB�
����W�À�\�{P�f�{�էչ�U�^�XIh%\[5��^G�|;unK�)8��ҕ�*���o8�?��@��+Z�CP4�i����"ѽ�~`�i:T�!7�k�T4&+2���3Ԅ�Uw2k������k"r�~v��^}B�	+0��҇�n���*P�ڊv@�V�ߧ$17���>\�_��T�c/z��QL��9����[	8�ڰ0�(��\R��nC��Ɂ�����.���9W����T�إ>�d�㜬�*D]^�pՄwt,إ�*0k���RGw.�n��׃%.��n[ݞ�,�� j,�6�D����GE��ݗ?a9�!N��:2���ʥ(g�-�Ha.Аʹk��T���3�Y����b8O�F,���D��[֐9qC%W��\��T��P�̂�Cl��巜�h�^z�sK��al��6��F�� ��"��2\�����+oD[�`�U�p�����)7��6T�O�V�pI3�)���·��י���=�{BD~�S��E�+� �b܈�b�s�^�qJL6AhI�.2Lj�'&���8�Ov����]v�(��v��#���<��H?��U�%eB�J�j4����yœB�1 �0����? T���Zt�+�����^}J>t5���٬	â�I��tj���Ĕ�DxXn�χ�V�j���R�>%����4^e�l�Y!��:Z���?������x!��8��D�PWt���uA�)X����W��jT���]�H宆 N�\<J�����璘���J�
K�㦶
�0��sL~ܲwt��?e%u�3�x�b����r�����Cy�{��=<�̅731b��r��AuˆK�2_`A����x�V�e�W���jK�}m���4<:b�K�s�9:�jU�l���s�H����v����ס'��Q�q!�ESjB�?+6�ݝI�CC�< '8%��)O��$]y)��R�.@�^ט[�+�u�E{F����o�ar��r%9{��B�<5�㤢G]<f��L��)�K�`����/�����ɊA�2�Dx�cl��d���f8�c��7��"�90�Hf��r����� �^dǶ��>�S^e������p����1I:'e�{ca��('�����4�+��E�C�Z�e e1��rg�c�=��6��((���,U �4���H��vi�_
�[���tՆө��uǬۤ#�mD�\�̻/�
�p��}%�<�6���l����Nb������~���?�<c�������Βm�+2;x��?�+�Dx��x[�uF6e�(v.;g����J�]�V0zn)Ռ���M���и��l	o���|����1��qNG�jZ�Gī��Rd�m@O��f=5e�-0���nz���h���K���������Ϻ�<�����%O�9��u�7-q���Cl�	����р��{}>%I�%�_�O���K��g���~T�z��.e�a��-F'@C��8�򳻿i���r,��P���h,[]�4�
봃�Sq����wh���?�H���>$4	���'r�i?9С�i����Ծ
Z9h%^x,L\���na]|�0�%Y��hꃔ�N�os��)�p��&;��L�9�����ɭG��|W&Q`D�9^�)gՈ�� +�82Ȃ�B�%�<%�
��c/����W��T^�:L�*�Ί�'�v���Ep)�:�vȉ69��E��a[
�6�\4{� �z��x$�o`!�r[�@_AG���,?��Av2��e	�ҋ�"ߣ��W[���#`ñ�C�%��R����!00E}�6KŎ�&댼�����z�B��`����z�������K�b\悗6&o4?k�yT��=�����]@�ҿ���cy*���$mϙ�@���׃�!E.���@B��K#�����l����Znf" ��RԄ1�"�H��#b�P�'��V���+��g�#o`����E)�����oy�_�Kki�bқz�RMI:��OЗ�z�G��4{���$�0~J�"HF��F��!R���.�
�d���o��,��ؙ|C!�VxY���mO1Z
�SM3ȵ�f�(Fs���$�����	�#T:��!�B>�:�OS*�8����`�"t�zZ"����#G���P]�[�uzQN�Mz{Y��^A�vp"�+=c[���V�;��>7²]�a	�#
O�q+!^��_%U�X�����գ$,����Wb���4Y���D7�e�S�?��il����d��#}�/(mW��);?#.��V�_-b��?+섚u+F�q��IO�T�Q�����E7a�`��R�Ί79A�g�F��h#q�����T� �o�@��Ql�=��}��ߚe�/��P�T�t�7��wa�^�˫cD|2E�U�5te��LXlxV16EB    fa00    20d09��D_�
ML�A��B\�����Z����^�xy����>Z"l�/���T��ϙ=s4t�#5���x-˚cv�cD8��nq��������k���braN�>N��7?|�v�$��ͭ�<b��0Ƴ*y�h�4ٌ��_�?Ќ��%Uz�k~�����b>��#�*ԞU�[O��:��s�'�Ŝe���z'$�}S܇' Z�r#���ՒX_Ȍ�J1��?�}��q�G3��67��Om�����Q��'�߳��I'��4�Y��I��F �Ox	�>�[�ա�2!�W?\�&��UR��ez�4s ���0^�U�_�?�Y��U��S��E�ؚ|ό��z������hf�_7����Õy��@���@��N����0��ڦ�:�CJP��J��e��)�S���?v@��Vh<���;���j@6~
Tg�G�v��W����[n�����_����) �����b,���n��6ʹ�8S�ľ�� XK �F��j9��0���>���4�����mc�4�B�z��R�������ɚ�>�Pl�i���uU��V�u�Qi�|�3I���y�6�dbj�Ӥ�<ZSzz-�$�r�h�wVJQ0E̃j�X�.^���o	O�����ke�n�]Q;�[�j$5�m��_K�{ځqdV�������P���+w�mT)���n�D��y��=�� ���%cs#⟇�Kt-M�2_�PbI�rJ���O�Ҕ�A��#P4#M�(P��q�*<m�Ꮥn"�g\���9��X�1
�(&Z|X~�=ҌT>]w�4����7l [Ԥ�?���T��)�����N��,q�?��:nQ�v� 6��Ï�:���nf ��-@�����~t{rs�ҎIR����è�%��yI��m����C�������)�F�g� ��x?M�C9��� |���v�$���>S�G�\(p��"W�v���x06[�����o3�*�����!��'�22�)�J&�o��Ϫ	4H��8A��'�_�|��"��=.��ߏ �.`�{��������&xP�q�n�Lu������@��K�]�Q:��j�y'i�z��r���@���#L	UKH�Ef��x���9�$4�6�d���x�EJ�'�ct�<5��ydnG�4�6`y*�	�zD�u5������KY��&۟�Mg��v�\�5f
�����k������ׄ��T�P��  �O���
��a�`���tD5QH�8&������g���{���sQ�����:�H-�4��<s[4%����5C�Fgh�e��DV�Ϋf�N�36!gF*�*���ʣ�%Y_��nZ�����A<�I�,���')�_1
Sk��=� {���E~)Uo���$�YhO�=X��3RWs[���b�	�*R���d\G�����J´�~*��t��xQۂ�
�^��Q���n$��uc(�s�=��Qd��S�R`��?�c��i�Q8��s���`�,��U��'*�7.����$��,���}a�"ߠͫ�^�w�v��_ �YQZ��-5�d��^)�fo������ee�,M���I	ᢸ;�mc�B�L�{|�<�V�I��Gj����.�� `�)��ݖ��C��l�H�������#�gLl�K�ڣe����S(�w�}Ck�6��V� ��~E0�o~�M͕�
S(�Ym��9N*�g��d ��PEE{��+��� N{����H�F�/Ҝ���ȇ��nW��{.�	��<������e��Ʀ�ӓ��L:��PW����X�脄��L5[�\ȡ7���ctM����N�;��=g�Ƈ(�Р�����>�q��^ /��o&�1��K���B[�,^�.즦�o�΅P�!�"�"Dmz*Q�ds�D^)�~���@�t���g���g@�T��WuR�B�u��ƁU�'i�kY�y5�l �/��꽚�Z�Py�*A?^ȁ�J��C���T�$�L���~���>�$%}Q�� yz� �Ћ��U:EX6�! 
oB��&��"�����!m'���e�!�C�Z�%���_8_N���mŃz��#<Q|�.�/�-]���xC�&��Ycנ��L�Ԍ�5�g��BW��C�ȡ>іw3��:M^�Ήa��eTs��nʤ�	i�ݰ)�3���L�ޜ��J(sZN��f
7�LѰ?���\k�3�΅`P~��z��WSO�|�*���PO��uR1P{H��Ǘ�Um����66�m���l�>�7[(�������~�T̙�_z���'�=S��t�ۄ<�S;w�A�Г3ɮ	 �bl~��4	���`HDم���+�f���ښ�����m�S���"�_��7���l1����;r�`���+����`����A�w�`n��z��|�n'P;����N���n���-�r�"إ{��0D�\8�_#���ܮh�4����m`��(!*�J�J��w��3�I�F�z�}�>��{	�����J�ݩ�ȼ�X鏔�0�
�z��FKp����qmc.����!��˥+��,�n(�D(�����9�@&k�LcDR����b��F��O�B*�A�Xu렆��סՊ%��F�/��d�`;E^�Xݦג�?�������J�Y	�����ȭ_�]�"��`gA����ER_��K3�s2Y���yT]d:v&�]�&~�`��n�����TZ��0Ŧ6���K�F#	J���'�O�|��|	�P���������G�$���`~�ǻ�>�o�*-I��$�������F?���4��q�O��&i���a�L����Ս�&w�� ��s��뱮F�?/�:���̫�m[��v"I�t���T�z�M���]���l��qY�c߀c���Ɖ�:�*A��¾�G��%C+-�p)���Pӧe�P��5�<�z�.s6+'�ZKˮ����̄fS� 9�F�\%���-�W���ځ�`�EWHlW�b"&�!{�A}�Q�Y�S5%����Vo��R���h6���� A���Xf�''Y�A�dl��tr��E[1�NG�a?&̿�\��7��c��,8�*YI]���QZ�N�h�.���m�gtJ�3�n�Q�$&��:�]��[t�ʿ�2�I�I�˜V,L��k�(��Ӭl�<�G�T ō����|��>��\g�$y8� 
)������Q� x��M԰����
�{�Y��fU %ilA�b)��J��]p0#�@{q�j����\���w�V��}s���~mN����a�q�n�_�m>[c��4�v��h2{��0�`�` � f+
;��d����� Rsa3(���\ɓ�@�99wo8 G�Z�TL��ժ�P��ɻ3B��V�]&�U��$���9��%�C)��͔4���/m�?�(nlT�R���������A՗�����&��"%���q����$�Yo�CH�g��_�[in��@��G�ò	�XaI'��5�c���o�RQ�O]� ~��M� ���<ď���ł���X�A�N?Ki	R��.ڥ>�w�h-��:l���.��@~ZQ���	����F�h��E �:�4�R�:n��[W�>c_-��y������X����fk����"�ZD�	�Xh�R�Du�,�r'� �/JA�����	� *>a��hǾ��ݟ�_�vAiI՟H�����No��f6�-Q�H~fx�$����;��3��̦�@X2��m,R���7�0���6�]��8�*����4r8����Y�O�@xE�0�D4{NP�����F��{�G�������6�*��J���xz˻s�kQ�5\��p��3�F5�}��Z�I�g E����si�H�6e�s/��<��<���	������`@��L�����\�Z'��1��!\��#}�f�{�K}���@ �+�ˑ����`b���8lF8�b�-Emp�az��G�`uƢ�%���Iz�'�{�#����*��4���;�{����
��S�P�����6у�ǆ�-�4B�3k�@���mʐ������ǁ�>o ���={��]�\���H����2g�q&1�
<�K"̀�����6(��7Z���xȠY>$����7��å��fp�1{.�6��r�gI�b�N�0	�$<p椵;��3�b��u��xpj��,�� l ���bn������t��;*���3k�����PI\������Re֫�B�8.&�0&@�����ƇK����R��p�6/Έ�fgOFG{��lx�u�?�I�|2���D׌!��elV�	K&9�)z�#bÀ"e� ����!}��d�Z��U��/o��%&:�u���7z�\6���
Ud<WSzZZNUo�B���}�g�<�n켕!��Q��.��>A-�}n7�>vu�!`	�z��m��q�h��D| �j��"綫������MU0lt��5�fp���?�h��M�mJGVfM���ycO��#	C_S�����8���:k�B)^+ὲP�_Q܂u������T�ҕ�_p�d6B��3�����}>�KmP��/{;~�h�V�>�-���	0p�]��!ǀ�g��l0�h��ײ�0�pTD:�k;{�|��TY2Ͻ��%,�g.k'զ�P4H�Hdpķ"�2���O6��N�Q��e�Ε2?�'�6P��4Cq.c*rB`,^�����;Nh�ዃ*���嚡ןS,������K�j��:�qb�_7P%\��~�A�ki�o`�y��C���6N����{�����zuOpQef:�>5�6=t��%zI�M�`�G� �2�ވ����B�E��������թ�)�V|��m�ن��|����eFp�X`+}p��=��$�sk�G)���l��>�g�=�>5ĥk$�cM�هVDV[�E7�mu�k�'�s�� .7����d���e�B:n�����{�Q�^>��G�0w�2��#����ȋ�IB���T� tSO�/��URb|IRC��mjH��@��e[7n�MfRh��}*|��r܍ډc�:�9��}\�2S�≑2pp��s�ubU�~N6.m����h ���p�%��fҜ�ȵ.'��`-�\�ZW���0u��H��Wdb%QEأU>����*��T&�aK�%dĨY ��q�t���c}5�k*�I�u�>�Sr����U�5h��ҧ[eH`������*WhS�a��	�l����@b��i2�|m7n��;W
ȉ���,��O�ޘ�6���wʦS�ZTB�U�4jԷow���/֙H
ꟻD�u�
0o�tʁD�z�
7}��t<�P>9���ql3��	��r\���s8���.x4���'�D�D|2N۹â�'<4�� a�����E�1���î��P?}�d,L���?����d��ޟ�>��]�x�����^e�nJ�(R�
�j�\�\��._�q)h�V>���;�Ľ�ﲎ� �sg�ҏ��T���`��fe#Gk��<���)���� �){��$!l�Y}����"̢���L
��,���ٟ�1 �]Q��A��ew+ A�m����~�4�����7���%z����[ň�%sg�1�2�4��I�����y5�kͮ, :]����߂�k�
1�댩%�i�uҤ�BϦ�ߖlB�v���l�2n_ ����7�o�:&��N$RT@n�kԆ���y�(��2�¢�)�!��+�d�Nʖt���&� ��'��,�1M�M����i�./;�>����4�V S�FqD"����vt�>zw��	 ��� xPU�5k���V�ꋜ��x8}V�N�0/ �����m�n�k� 3��$C@��������\�&|ی�lC�e�Oގ�@n����������,�����J�=�߾�t�����u��W|��	�������J����h�fFћ3��Yc�	�����Q�k�n�a��#!p����l�?v�O�V7�g��4�f���� �^����xE_������ӎ�]�Z�I��V�����Z �Y�~](۫�d��d��hs,�=�C��D>��ROK|��q��͘W(xf,e�-3P�|a�!���a	��H�٠½jE�:���Tn+����ZH/�t.���J�Y�4�:��M$��&ڊ�W�u{+�i?᜿��?r9^�ݑ����v�"�֬S�\�o���d��.��|�U�O0|��v�ӄ�ѭ�}og�ICfA�<���� ��7[�[�l۞�w���~��Wn�9�����6���㓷	�h���m�K�e������C|� ��M��=���
(��ݸ�ճ`��G�\H,���i|�P��-5��������Da׾%�B*�h�>�b�y��̆d��@�D w�V ݥM*����+���֖��!����o����n���N���"�(w^څ
�-�U󶬘[M��/G���s�h"��%�9x�$I����a���B�S�j!-�ËT�9U26ݻ��(���%M�`� ��{���r��X�����l�;���%i�����3��I������:C2փ/���L%h����ԍ�'�3#�-����"R�^<�wG�v"��r4�@e���␊]�s�/�{��C^b�_����	�#'�徛�kn?+�̣+��k	��	&���	��n��SF�s�����>pw���k���Y���_��w�^�b"��|�R�G~�>0b|͐ʆ�ZU�/4�IG;B��E��Pg��W��@�êy���o�5�h�U!>�E�!$l�${^��x~^?�fH['�(�rN�o8�v�6)���XC[��'i'/(9�>1�kMo]���[]�^C e_��ur+��&��m�$��U��y���N��3�XؓО�6o�]�]�i}�?֣y"��W�y�Q��=+�O���X���M����taɌ"�?tȕ�#wÛ�;#�G5䁺�n�̳�e9���t�7�N��K��3h�[���҅��rP=:|�c�CG�⊭X�C�4�����B]Bx��K�NI�T��$�S�#���ي��ȷG�t��oRm�"}LO)j�χ8%�ގ���O�\SJ%p.ƿ��<��9`@��w��w�#��t�#�О�NTFڿ �~}m�e3Dx��K�(ہE�#��#���hY�CRJ��I0 dr0���#2�n�S�(�k_��;0�ݡň�t�`�,�T��D<h�����
� l��sn������om���V�*�#���5���U$�q���K���/N������ ���k���F����}s�׌�,��`c|���E�Z���ٲ�O�2!
�)rx������C��ȢؿҕZ�Q��:�e��X1��^X�d�'R�,��S7����F뚶t)�'|	�8x�j/��Ə��$�_���	��3i�(�84�N�������9-�	�[�/G��,�p���L  �q�&���[������e�\�7��I���+f��܎���0~h}��1$�Ǻ[�ɦjWFy�Y��sk�|�9�W�?���)��:IڧN#�����T�\Bz��9���d/�i�s�s�����$M�j:߲� �F?Ɲ1ɣ�s�2�^7�,����w;�{��:�L��V|m	XS�O�x����lbp�xD�z~���2�=UB��ڦL�һ��,��x�*ĠH@)�.Y�.c*j`�� ��-���Gd���bg&�������Nd���t�`W�r����@"ؘ ��ꡥ�w�����o�����yX!/a2>x���H�b3�T�8�1�����vl!�'+ñ���#���.q8�5���Yqf�����gA���ޥ��j&�����[}T���x/��D�8�_Hvl���#��	|��D�c?�N�9^\�~�Ɓ�r�9&ѓ�ᕒ���G��d��`�@��o]9�<N%���_r�Ď}!]�]B�ߘ�X�`��_;�,�^ҵ��e�x�)���A����k�v����j���Y*�kM��6��e�z^�m��l�J�8�4��[��6^���@�����ڹ���G�th��� 88��[�<�̡2:Hsl�>�B!0u�����%����s97�p�v���Շ�%��v^���G�ϪL�Ds�j�N�y��2yV�)dPR��-�cSg����\�BR���?	#lbzOߑ�����Z���{z�3x�n��|wm�XlxV16EB    fa00    2050�k!��ۻ��4�3f�Ȧ��`X�w���rmUB��� �wY�� =ŭ��أ��SĴE�z�p͗,P�ĝ��(*\&�6��nl�=$��*�zg(l���o�o���:�6�UTL��E&s����%CDJ!I��kO>��� ַ~u��P�}6x�\g�.!c�<k�oN.��!�p:>1����$�k�7:^.A*��,s�Z����RP�w	v�w�9ήM���5R&�Ip��4R�7����+�G]�m�K]6��A:�|��\�w�����O��/�G��.����hZ��x���O��9�M���r:b5 H���:��� ��9��<v�������By���/f�eeɶ�����V���V��d@���kR����s�jʛ����5ы��3\��?�F�4����n����RFh��Bz�G�h���-�"��K�_ܱ�kr8r��^��ēå��|�Ӛ?)+"��|�+.7�T�J�\���o�@�t�w��o|v�<��e��5XF~�ak$�7Z6�'nJeM\m�S(����N(5��)��ݖ�TyA��t=���<Y�l���?z�k�hO"φ�OT���5��1�ҫ������lz�	��Ul��z�Mp�_J�o-ڋ'��Y3����<�[/���R�l{�x;��vo�b|�j�w��c\�e� f����f^��O��b���&��;�o�{���  �u_�-a�����]������,<
D����ԥ|��M,�����c��2-�I�Z7���N}gpm�lg�f��1�o��ʖ�&��P�iF-���+�/��&̙�?�+Ŗ��I�ƽN\s.戋��^�k��� :��F��	�6Ld+�>޽�ܗ��6V)�7�`���d��Y�PӌQ��p�HJ�N�S,���'��%fOݫU��\��\as�7��gl��2��7b����KX-�1��hV[����}�(oo��;!�PP�g�����N:�m
����F�nt������f0�CMص]���2��m�^�Z�ʹ�&%	��W�^u"�xቚ5*�����jK����iK��4��K[���c{�B�V�@<>�Ƿ*�n�yq�l���¾�4z�B��!���_����vH0<�@�l�E�V�
+v`���f!�h/^�H��'�	 0tG% «��<*�l���u&Ơn��BZ|O�v��4�m�θ���&[vJh)$�t�wdpʣ�ܜ��i�Gm�)Xl;?A�8�7*�f|����w�r#=qfdn=�>�Nɘ9c�+�z���M��h`���}g`�n�����S+o�C��&)wS!J�|C�~������W����5dR����٧*s��˫���,���.�T	��f��.M p� E<�U��0nf��Y+"\cY�ʧ��K�*���`hs�9ͦ����ŷ�_a��4�	v�m U��G��\}���A���ra`:�ͺ���m�b�kK��S����o 4�˫G3�[�s���ɜ/����flA���e�C�?7�? ���t\DVb�4��������ܥ������� ���Y��>&�C�������q�
�% 9P�͋C�	��w&v��#�ߊc�����u{R�� g'��ԁ�G�e'��B�	m	��y.wΑ��g�KF|��~4����/uX�|��U�RW���j����Ɠ��b2�*q>�!j��>!��
Km��	HZ��Hst
s�:���6kDy����5b�z�5>E�@���M�1<^�P��F��A�5[ݰq�8�M�%.6'�HH'�'��~sQ<�=Pip�E5 o�c�&dя���siF����/5k�g�5���|�G���)�
�X%&��U\dN�mB�EV_���0��	�)[�h�k8�Ҋ����x���ӕ�5��^�3#`%"��G@I��9�d��<�Ru�dS�x�A��Nz��)H&kӫ���|�c�⤧R�S����G�^q�� '����I���t�+/%-�=��Z��z�����˒��D�}�8�T�Wy<C�㕡$�~�6/T_�݇�l���!/lT˶�<(`�"�G�#^����R�e����7z�ucǬh�;`C���T�%�uF+G����0����3e��J�W0]O����$�v@�#�m|���JۖS(K;�Kp�Mq_�@�͆���*x� �D�H���Y�&���*�/�tr-�ad��hxz
�h���	`�l�)y��Y�SI�cYk��qy��"{H$�x���聮�-!*�,���>�����Q˪�nR�>Ÿ�,�9���w/J7m��!�̮��l��S�[�P�;aM�5]�cLU���̍�Y��`�&�$��'2:�Y��V�.{�J��nc�8ڻw J�n�3����Ї�s$��i�l�c��%��k`69Nw�KT6{�؟T������'�g�!@yy���'�9�0�hp���P4ϰ��W3�Yx9�[p*��hxI�"�>A�u<79'k�^�Vr��$-Ӗ�wBZ.;-*R粎��Go3���K̤^v�� �e�WM �&q�'�df�WI9�v��HE���xP(A�"�3$��:t\�M���,�@+S��,�d�G��l?x�ʼRq�"�����@I  \k���543�����{Azj�œ��VD���� 01t���,�Ib��E��+}u��,� ��$��S����uny�[�J�F]'��y�{z �]3-�fZ�C����+a1±l�$bZ�/x�7Y��L�Y��[ʀ�;�:-0w0�UU7�px{�N�:��� ��7��2GP�R;V���	��lJ�;H��g�(�6�Vc.Ʉ@f���:�j���5щ Mޤ�@,�ـkO3FӃ��g���a��hm��۽7ϝؽ4����W� e��P1아o��/5�A�<�'N�i���0l�|���M���0�"~�y�&5��I��C�s�x�]I�+��T��`f-HdL�M �o֌u��T2͈w���Һdc���A-���Z�y��gm'�)�NR�3hg�S�����;UjY����2���ԟ;62���GLޱ�$+�M�|�2��H�(�>�L�z�6˲q(QAC����C����r�W^N�Y1� �-��a���2 ���Oo��!c?�y��h�L��}��Hn��� "殆`�0YG��)Kq������ =�Rxj홰���s�-��cZ��'�!���sנ��#��B�G#�}�]T*_�������b��;詔�'W��S��Y�$���U�����\���)��>�¼�����25���9��p�)߮[K���f�5��N"�c5I�v{��\��l��.�c�v����V0ladxD�)��"`����c#'l�t���AH���ڪ{϶u��@#�۸e�#֛��K<��!�C�a�H���4*p!�C`�Y����D���4�&�(��?��UU����<�:~�c�?�b��� N߲�XykFr�������{�lyEM>�մ+��q[d~�#�6m�T�zܣ�����a s�W-<V4�Q�psJ�uo���AD0�7dSO����p#x�,-�JQ���V;6������ZC�ɵ���-M��G/�1C���u��eP6�4*�K���~��İk��[�^��{���j��=2%��Y�����f�F������e�;B�h	9_�������lh~��J@���/0�C坺��ڃ&��;�d�M��`c�L��� ��(��L
k�X�q�e������9��yv&}����( �,��`ôqJ�Y�!
��d%�N�ԙ)�H�nHN�W l��@ldo7�1���Z��49�H�K��;���7��L|�h'gaE&ZC�.�z~�����}r�C��~����tK���C�1�-zt��O�eD[����ڢ�������s<����p74u2��:F��W�e�3g�S`�K4�N�u��՗ݰ'��[��)��C[���^���nK;w�6���@)|��b���|=�/w��xb1^��2�K�������4��7G�3!ӈmb���֊mh$�T����܎]B�A��õ:�s��+hbLp�ESz���O�x*�b�M�+ov-z8;pJ��r?:�y�?�ף�R*�J���vBϱ�E�������I̖�L��$>8�i�w�&��B��@���>isV�?�g��0���5�JNb��D~��	mfr�����Ae�7	�N�Z�=�Nz^!��g���!�g�ѵ&`����g\c@b�������հV]Ԁ�irF���Ԡ����CTT��$�qw�]�H�X�x�>�ͪ�$���X���X�Q!���`
���9�ؙK�X�08��!TY�P��x�D��������RP�*h�^E (q��H�����N�@�������ˬ1B/��.�����5����zT8q�+����>��bV�cj��B<W{="7�IO!����
�gY;|49�hF�Ũ.��gY��㳰!�G�v=�<Y�|kG�K-�a��Q߼�}��E����aO��'X���,�s�I�PO�Os�0��;�CHp<̈́Opa����Ƴ���A@^�7����m�����%���]�=fDO� S�]9D@��P�dS�7;�;!�^͙|z_�j�Z!^A��Ͷ�-�c�/4qZR����|W��at���	��LM�b��xeq�A9��'�8�K�(�-M��ԕ���[���u�\�Lu�C���m�t󡈡�<�&b�.x�?��4]
W���b�Q�y��Ȱ-W(D�?���j%~ l<��5{�����W6�"X����LU��"���ݠbM>�v^t�z�d�Ǒ^�5ŵԜ��M��."_O���%� ��z<e���n@2�鋺 �Z`���v�6#8&O�{�R{ ���0�t���_���B��	wք0Rה��;�%��ڜ�Ъ::���a=��ݦ�N}���;��5�}����R1%�DWϥ�%�ll�X/`6;��v�ȧ<�w�����V(��A�\���D�������~��1���G�<��r�WVz�:*�̽��Ji�&��|`3��8���4��֤�ش�
���KF���<uE8����r��R���e9�H�J����w*��x;K�K����l�$W�F��x=<�%�VyF;9k�m�^��R�!�����=�9��M�qF�lI����^��iUA�w�J[�\v���!��ֶ'�tZs���ʚ8򐾔\b?�W[��U�=nX4�����X�k��e'[�e�s�,Ĕ�j�f��#����?����]OQ���1�{���,^���v�����b6 i.��)��׾rAYu�`��������Zrm�^��nW��4b�����Q���:��nX���sI�:e;�k���F�-i0�%�p��-d��!�b%�>ӏC������	���?e����0a���Bu@ a<~=$欉��z���,>V1�*I�Bw�p�NU}F-�1UU���D��QXn�H�E
�Yf��xb�C4{�D�/]sY�v���{���E����@�� ���P��gZ+�N��羃,w���rl4�=���'84�a���S�ـkcp<|��xQ�+�l��^�PSVJ�����?����k�YV����}F� E�Y��* �.�%�UF��(@���[(�$u��ß���X��*�����)쎛_�Odv���lA�	}/�=JN�܋����ƀ4�1���掬o��9>�I;�z�qT{���"+� S/'3�H����=�xǡm�/U�k��Z��O(��-"������Y�� nh:!vu{��L�~<�*��_:���!��bN�QN@�)?��yb������h�q`�
r��U�w!�a��U�0#�w
Ѹ\;��_8p��ll��L� #5���Q�4ZS��rTW_0�S��7�ZN�Vee�ȍ5gq^���Q�k=���yBE�
���Se�K���i���K~"R�AJat��e��⽩��`����5CQY��XH6����|z���Vy��)��I�e����K�ϝ��-�{?�)o��l�p��]���7%��%�'����z�<�V镡��������G�-
��4����>%� ''B4|�T�Z}Yʫ��
��t��w�!��\��]n*UT�p��U�O�CG�v�Q��&�z�TT�1�m�`���7$��5��"9O]$�	OXl͝�e5����'�=k���q57١��9�;$7�i+����
tqk�r�������[}���Ʈyp��W���<9�@�^AUswA$��^H����l��݀�Q"]w�"mLc������KL <=���RBp�7���T�#ԩ�����ȧ��;���Y.����Qy4�o��������pŕ�]��b T'�
Y�[��Ļ�X3����l�}��S�x��õk>���l��Ch����/V���3�0ַtJ��u��W��͵=j��N�r���xC��k;Vw��ӊ,4��'�K��O���>�Op����ft�lo�3��j���L�KS�`��\���(�j�S� 1[A���2�u[\�B^�@$�M�Ol��E$f���0�Ϥ�܅4�l$�E�����zR0I���;�*������^ FX�[B�ou;��m��VLgtk<�^�j�ט?�~���p���f'���Ɍ������r�}��Mk�tKPWq2���߽B>�v�9�E(BĜ���e���� 1`[avKpM?&�91J��N_�s�&_����]e�,]��=2V��Hs�%32lJ�S8-\�<�7���_�И:Ѷ�/Fp��*�T�us�=� �]�8a��pPð�
�-��h�l����7����"
�N8v�5?GI'W���F�D��gt�� �$�� J6���0ʰR�$��Snh��*�[SS� ���8@�ׇ���QU���p��/fa���O�I�S�͈.-H1Q�+�^��^�tсt�dV��r�sk��q�dL�L ���+F$
������������P��n�tC�1?��7�s�E����I�����q=*N�V񥨎��b�j�Ǒ�U9�p�ɩ�=�w.���Uo"6���eM0���~�� 1'��W3�
����\���D�����m�a<B=J��"��;f�R��i� そ����#���ZǫF?l�
�u`TD��n��BA׳�߬��}|��MN��Wr�rk&���YL̲�Oٿ��z�HC.j��BT�T�>z��E�!�\곊������;��7	����bIKC�8Bdy��ˤ���+{��hjF�%�x:�iE`>Q&L�:ln��Ӡ���b���a:��Ҧ�a�rz�3�1�Ѯ�|��rK����3,�[C1:�[�i��1����=̯ʂ����@P[a���
/2U�;1�
H�8�q�[�ew��*��t�Q{>�o�,x��p�^���W8�l��X����E�B�#���5�ng�P�`/��^�0~,
���� �r�����6�ӧ��r@�̲����1n�3̇!�׹/p�V��˲X����G������w/��S]��z��H�/�"Ωl/����o�:��������@bܝ��H�iƨ����� /ŝ���Y�^E��OvW�t���ޏ�kf�/�^^��s�D�G��s!H០X�{�+�o�k��z>�_d���ٓ�����F�{1,pN)g�f��P�6T��5�q<����f;-���"��ki���?��$\��J�+��;O(pt-$�	S���7$�>ߊ���U���KK8���_�cX{wR����z*��4�H#BN�i;I&�KH��,�Gi<<_cz��H��c�2��`��d@dz;y9��ӀZؙ�I��UK�w��&�m�X�M���c�>�pnz`����r��Y�WT֧,�b��1d�(������kJ�ht��Kx�b�����C�<�s�62�u�ͦ�{l:�UF�7�Ee֘���J��A�ݍ��[��i��oJT���RcG�2
���rn�4r
� q�Q�1�&���/e����=	o��b�6 �j��oL�ߓmc�Щ�54��XlxV16EB    fa00    2120��������OZ���\ac^��'U
b�M�;�\Z%d�$��Yt$>��K�פ
�7u�9��i��7f&���-��d�.
�%�ɍ�ۜy�'�w�����ܝ~
"��bɢv�ګ��_9����)	�2�,��>-[�:r^N3o����׌>�
�0�>���G�������*�Z�T��UW�Tj1�A+@���G�s�:f�W�ŵd��\�=h�5%�47A_�	�=��G!\l#E��tWC���:2ޕs%r����]�7��MǇ�ݢ�A��U.쥦�C�V"��ʩ%�1C��s+0�jPZ�A�G9x����C�!,A�п�mN�����4��ԅ먊�U+s%�5T��C�%��}7k�	��$����/'��f>�k䂐oQ{�z��7nUe�z
>��^˙�c�4cF0�҅бdRKs�� ����&��\h���>�'�H�' -���${�㞷���cJ�2F�>�ᝃ�"����OƜ��Q�G5񔠯(f��2�L`ppQ�abD�̘����i�E�����dZơ���F�ٟ�xxJ�=r�ŖdAY��=�W�p�ӓ�c�e�LI�0������.u=��L/c�D�c�eZ0���5|Q|Ϸ�5�_<އ�:=��!��!VP"["H���xZ�ڄo_�کp�}��h~J'�\g"(��Ф��P�7C%�u&�|`Ӳ5����`�m�Qɔ9��E��y�4ꕼf$��Ϙ�W�ƊJ#7�{8in���~*҆R�����V�)H1U:��DI�M�6z�R�h� �C���ʴ�<�^������P�o�E��-sB�(��d<;e��S�1Qt�(p,�!�,W��g�(C�r�����g��0Տ։���� �*�B�>�1�ʤjkoLBV"%���B]a{8@C�>�����!��hT��$c]���;���<'ɽ�U����{��i��o*17.[������5k�����[�(>�҉�^�?8*#�=s���K�[v�R�1��r����q��9,>Z=_nEs/UI2�p�>��K��1���Ĩ9�@eXE�|a-]���c����T8I>���Q�P��G����V��#�uE�V����(�Yv���<��~(�q�t�,�6�O%�H���"1I��D�_+��煝�o+|�c��q=/��õ�p���X�M;�	��R�Vu�xR�g��i��Й�+����8���&�|r�� ����L�r$ cB�c�Zd�َ�Ӳ�a�S�a�������~��P����H��d� 
r�V{��8^�f�Z�4�-nu������*��s�- �ۢ��qZ���H<�
�}���J_�U�K_ X�kTe@c�I^Um�Pھ������~h�A��pby��ixLj)i�w����p#���2�??�t��W7+�s\�I3!��f�ܩu,�З�Oh%Y���~Cp��-'V�³= d���
-p��=��uP�KK\����w��y"�U�I�~�T'ճ�+����-<U����E;�w�Ԫ����]���w ��fB���`�燛�%�}]��a̱�9�mx��Qȅu���;SLTՀ0d��G�כ�pg�&Qi�2`��r�If�8
�t=#=����!��DԬ�|{��;=�q;^��-�/����;j3��y���9��D�<�\��^�"%���l���bl��L�ֵg��E�eK���D:�3��J���X�P���7�@Ʊ�f�e��Ո�׎��q<t`^��MIbEzGu�Uvl@��D%��h���?�Tz���RJ�TZ�1��dr��N�=�Xb���8UO���J1�1b��O��O��Z��[B������3�*�z��q5
��M�p+��6�1a�=_K_����l*)��ύcۡs��t35]�u���Xi�&J���� c� �}�F3Ƹ<���h0��o$�2C�U0���|�0�wV���b���l�:�� �;�����|b�4�M��D�&L��}��H�$V��_P��K�����I�`15eS�1 '
�����F`@��ʀh0#J��*HG��Ӥ���on�Ih����/� <��z�c����>���.7�Sқ6S�����P���JHVK�PÜ4�Rp�;��j�#_⤆b���Jx����m�5i���-D�s{i�H���TI�`8#�{����2]O�7�
B\�v��8^h�S髠ێ`!�|/�U��@�;Lz|��/f�]n�/QpTϡ�TX��_��|q�ʩ��2��!C&��㐣�M/�z6��; ��xg�9ȓL��=�(�|ʭP�,��W��&����d�J�-�,�@�Y�Bac�V�5H��x���X��aL%Y�0k��B�����������ʲ^?U�2��6�1!1��ݘ/j��� ��.�T�2�,LΜ@��G����TM��y�/i/�}R�maY��S.�����`p��7��jC�X-�,	�4��|-a���>�T��H�两e%���P�	�����M+�a�
j��h�l��k������Ğ�<!ib�X��<���*�
;��z�Z��O-{�[�8S�]&��U��x��	�����%)y�r��HW���о�E���ᖒJ�yEDEb���e��k�#ecZ�R�UHWQE�!K��JU��ĝ��X�Z԰^�^��؏g�8��R;-����<V'iO��X.Ͻ�[p��g*���v�bg&��
D���κ8��0�a�2"w�ݽ����1R��nw���Ұ� 'm��ں�9r	1�n!����X+ ��p��Ow3L�?|Z"s��.u�PPJs�_߷�9�BS��{�Qִ��'̌��$M��z�dB�1r�|$���[/��@^��=�<|�WI��3	�4	�a�ޟr	 *vxU�|*$��UN���'T�����o�k�	[�؟t��C��i�M�A����L��Yb�����
����Q��
=���m��V�i����oP��q�*�'�pp:Jb,e!\1������� E��ԩLq�3t��cLo1��ѡœi����A���U�ﻅ���4}k)ԪYg�F�5�([ٸ�b7�u��?{��H�o�ӭʜ6J��@}~<���aٓ���WM�l��#��� �.1A`X�_������4�+F���?��%�,I��ȝb΅�{$ň�Rʐ?�!�[u�ZM^�m�h,[n�~І!]%�Hi��Zeܣ,V߁���̝��j�����l~rV�;�	H+|;Ph�k�
`[v�������9R(|5�,�2�n1�R����������a���XtR^s�f��.���2�e�'��S�b��-g�Kkܓ���)�ȟP�-���;Ҟ�Ι�*2t���rc�%~��_�i0��$�X����%A�0j�o�(=IX{�m�8����.�˺g3����%�, z��Hw"_�hq�sf�b�VΙ���#�6_k�4J�a? Y�KF�5eyІ�N����T�q�]����WѱVx��߰F쌘lW��)jGbkYޯ�\�Z�3r��)f���}������,U�~��9`Xy�E� �<Ⱦ�Sj��C�v�TՄ�+S=r�(!a��,�#V�Ӵ���I
=.��D�.�pu�ǀ��J7ć�(��V"`��i�����y�4�	AU!2+:oi��B�
�^;4�B�8(��4R`p̘W��J��P[/�R��d��|���.Bq+'$<�clu	�J3d�b��a�����˖8����/�Lm`
1y[�g���axn�$���֤�d-�Zc���?4��k�˔�w!_��>�pDWj���)�L��!]R�&x��B�K�z��d�zvx�I��~7A�~�$z�Bc)�?���lb5�op��<��x�a��ğ(�M���yY��l�(�/�y��خF��̺KaQGuThM� 3�\U��C���3�hh܅���d�h,×�����V�"��P��,0<��:��4m�/���Gk��_�%����E�����
�Ie@+��=�������^v �c�W{A��,�����Ylֲ2s~	���v���<DH�4�����̊�5.D����qbガl�T3鍂�2f�����%
a}�W2o���Ϊh�!�Gf1�g��6q�������K\A�h�l|���*��(	h�̀$�M݉� ��Ќ����x#v�����,w���H�9%+௞%���I
k�c��r����Y+�Z�d�b|�}~�w+=Z��ؑFN�m�%Q��/bp���o��H�_D�Rm)��oR!�u[M���v�1���Hw9~��e#�
�I�����&b��%��:��r���~v�9J;��x����*�Z&~-�S�5��մ�[�n�yqU�!!{��V��"?�5�����
�w7WJ]97g����mW�>#�{��O��v�-���?#<	>\RE��
H\p���,��=a!A0�kF(LBN�H�/�yN��,<�*�nC��<�ў���I����Cx3Y��p�ݑ/��uX5�gL-�]m�N`��0�������R�1�~��q�2�L���V�	�H��
[/ﻙ1��n|���<�|��P����'qny��B'K���@\�f�+�{|��b�<H��7����1�ij"�]i']��c<�U���4��@2"�X�e1�[T�+>���6��I���4N�9���t����T$��3�>G�o!}�-����J�#�%��Cx�{[k��3{'#�<u�CHQ6�\e��yש|#�jQ �b��"q�Ax�=�6�'�.�'|���R}�X���w���(�L�܃�W���-��sy��lpq�f�!VJ�MȲqH�U`���؉PX�L�k�s�E�â~��2�h��2�ܾ΍̥V��z4�x'*�=�(���ĝpYC�a��W�=D�To�@��t�	6X������4'pi��0��{��}F���+o*K�����+���*<T��;Rs�v�cc�|�q�^²�[��u!g}�C��>����1�=E
��!T��c1.�I��|���h���V{��u�4Ldc��=�Ј��b��*K�<u�.��m�(�� �6\����!�����f�t/ p�Zi���q�$g.�ak�6»4�'
��#�<���������VH�I�O��UY�vr]Y)�1���gKGdQ�j�c�zP��P�A��$T��F"M��V�+Hy�p�
X�ކ�M��-�~�:@@�끬y`!F�]ְ�93�~�ydh*a�t�!��]���+�����#��+����8D �	�B�	 �bR_�����\5�\f���M�~�&;��:M6/�l+���1Z3�;΂��h0^�Xz�f*>�s"4IC`��j�k�pP5~z�7��x�	�8̈ �	��-'�Xߕ�YD�h|��h4ų�^~���Kք�w��p�C�̓�TO6sቪv3ty<���>�N�Y�c/3����8V�wH���%����/��(s����g�����z�����~��QR�f#�q�Fy�ːa�D�WCy��_ ��\���W�Fu$0�J���^�5<r:�K����Oҝ17��B1�Sj2kٞT7�@J~��D�SA9�dB5ƕ��m1����n�;�JNЂ���e`�fá��Qn��Qͦ���6��ϥfיG�~��z�m\�jM̢��tC�8"W�)�m�n�ʸ+ḣ�vu�w
�8�-����?�A6�o`��?�9���*{>�3��Oin��.�Η���b'(�{�X�{�����zPlG+(�/�$%�I�Q��!�
��1m��8���	}��v�
K��A�݇V}��e~$H�hYO���&�����o�C�yZ[+-��F��IGя"[�>�.'8���p��;�f*�M�7'�9�6#�3)�z�]�Kn��"��99����9���ߡ=��7e�s�u�3+ :�F�,;/�I�@�X�s�D/OQ���f�u@�@a�H�� �
�<��	O�U�F��y!�Ɀ@�.�%�ŝ,�ok-O�n�/��6�΁v��o�55�æME�3��"(�[�`&Av����G^��c���y���A}}44L3�%�^�K�{š�3�����$(oG��t����S���1�$���i3*�����SO��=�6+�,b�*���z<ޝ���vhq���z�^��t��!��]��{}�����o�D5��
��8zYQ�j����k��O�����V[�x��v;�H�71c��H'�ǎ���*�Q/cV��Ϭ�O���w%�7�H�-L�<��&��Ia����d��p+*�+S^ j��W�l�%kf� ����Ҷ�Gƭn��!�|��8)�Mz3���!d�fR��1���y�-������ׁh���4ռ��_<HT1]U�&�7g;�m�����7� �D�GT���]���p����|vG\&:�Y$j��}<)�wW	I���:�<n��XI�`^����F���ʲ\� )5^-��5��ʉ���5f�7���H�ɼ*X� ��mjr�$��,�[��2C�Z9���ËS&�и�ڣ��A�?-�%H����7�^���_TG�#4icd�6V
]�����ʺvA���r����\T{��r\���*��� ��J�tW�:���p"^�J*�z�ė����K.�Ǒ8��Z�$���9'�(a�d}0K׍Q��(%/�S{r6����.�)����C�D���0R��M_����}�Zw�(b�p�H�8 Y��c��X=�A�/�Dܟ�F�`���Q)��K_^��T����zT#�����g���gx�To8�M+-���ז;J7�튚WAM"k!R{���Sp�)ºh���(�/?�4��j�瑛�ё``B�=j�1���:��LGT�We �l�l
� �nӦ�VNZ�� vDR̊I͍x��B���{�v7ȂH����L�L �f���h��8T"��,Z���Ŀ�r��)��ϗ�_���(t������tX�A���|y��Z~�u̞>���0��{��ϛ�E��(A`~�M��u3��۲<��*Ή,��B_$"����Uc�#x�O���
��AJ�n/��ϊ�牥?�%��dݫ���V�U�@Ԓ�g�A��:g���;�)�(q�̈jB�e�l��[��~in����DŴf�M~��OF>�G�rB������k�/d���m� �Br�H̐%e�̵; �6�(a�!*�WzGe#�(5ZRla�}p뿽��pֈS�]D�@�cݫֈ}J�mS�ɪ4|x�?~oM���9��	��q���I����8�<n�Og��K?�*�ŀ��Q�"d��b,l��te	e�����anc���k=�4�@������,+n�Ecn'>��/���3<�pr.��%�I��z�2�n7��g�p�Vz#<��1N��r���*�@*�>a/��oAMa�aJ��HQ�Ʋ.w��v�@~��#�\�\�%�[ܧ��/~Ǳ��vDռ�&�� ��g3|�"ّ���&,p6/	�\׸�S����g�f�Oys���T�m�c�Z���u�Sv�S'��.�U^i�&�(UVH+���R@����zq�ڻ��4\�*<�j0|�顤�Wy���]q�"[��e� �-Z�� {v_��mY�;�{��UYB��x�5�������r�R�f�x楤ո����%�V�p �[�$�M���58 ��jI�ܔ�2Ȃ�����l9Zɨ�Ml��:�H� qN8˗b�7M�s��uN3�C]'KvB�2�� x��䌕�C�7G�QIH��Q��h�զ�U�,��C�)�Vm���	�72�&�5��֩q�O��fu�YmІ��b18]���+�sY���r2� ��G����VؕR��Ӈ���Y;�RSjf�B�njN+?�t�5�T��$�ި S+���h
=V9�������^ �5�'8A�j��s�Pnm�b�^c��l�e{���(Z��S}e���,�w���e�%q�o7S���]�ɇ���[4;6�2����������?-)��U�ځ!�0:�����rW]=�L/s_\AړM�`cm�[�r�[j@����f*�#,蛦$��u�����j�$R�㤶���o��x��R��%�(95>c����Vm�����E���h��7�X&o�(uy�pUt���1��y�h�j��tdyX_�����lP���G�!j���Z�Q���ɶE�#a�x�٨�J|�k�Q V\r��Z����"�EB��W�[Z'|�þ+�GnJ��9~�74Wɛ��u�1%���ne����5�W9�a`u�c�~����,f�e�&�G��H7V��a��2AD� d�XlxV16EB    fa00    1a60�N�81H�E�20ӽ��f�T��uK�}��v����z%R�tB�E��q�lb!*���2W^P�v�al}����=Lx�j���b��d��̌��I)0`�&��n��F#f�
-�Ф`�|�8/^�XTy�gw�yq\_�y�����*����� �Ύ��<���q�vQK�N75���e�6͌bI��.��!�!��\�FR�e�"Kq����z�J��1L�����ˆ��
)�~�yM�Y�`�S�h8]0��^�n�(yC'H���3�A���f�}坡��e�﷛�l<���י�7cOp���v:(��]���;/�l�v$��s��B��Π�F�U����,0�п*2p}�Pk�
����h)1�9e�Bͻw�,�0ܼ�o���^7j�n���Q�4�5Y���=���W6:ښ~�0�V3�ft�ɳ�oZ�3�y#(8��������nS+�S6b"��'�~����+HM�8�q�lj}6�[�v�ı���Y��*DU9ԫ�?�9Q���.�Q�|�&���43䆴���%bk-?�
:����j<� �Q��Ч�ۑ��)�P*"�hY^N�Mj��/�X��J�����*�VE�*��'̴��u���]�|�
A'Ď�ʹ�7-F�bٲŎ��()M"6��$=xbת�ņ�I���C{̈�>[��{�q�M��c�r�,�\H������^(�d��3�9:'
��9��u�5�Ԝ��Q�R�6��"�d��L�#�RkN�@�t�E�rB��OZ#�(�#&���gY��K�y�\k�P�*�Ώ+���ά.��Վ;���{��匸����P0����@�d�9���O*�l�>J`e�p!-g�"�BvB�RA?��K�ƭ�M��˟�(��cY��/4*M�O�O
	ᩓ�#
 �DM�խ����a����݌�_H�轇~����oT-�jj��9��́$�t]%��RJ�D�M_!�1���mbV������g3Y��̜��N����ӔVY�g�m���z�d[{��438�BI������,�f��RέZA��Xq4���
@p��H&��ut	}|g��"2U�K;��39X���D++B.�:�a"���] 5`�b��N�񊠵Hy_T�nݶ22BP��0"Z޳Cj�ׁ����%�/}��$أı2-w��ra�W�����Kt?��.v4��g:�Y�k�5���4�6���d[��Z��� ˁ�g+\�FVDa�)�9���e�RD����V^�P>�|Qv�p�ך*@2
����<F�Y�����~&�ņ��*P-��'PİM�����!�������m!�C��(�X=���
���:���c	�8�#U!�`�SSȞ'��|�M�Ѱ�D#�9R�V���0��E��&	ڒ�,<�me��4%��'�0칷Z�wِ�{
f�!+�I�.saUd�_���}�8yFM�/F�[z�kT+�k�.f��0�oj���[e���;tAb�QTT!�f�@��Ģ������5��@�c���ӛ�a�ߛ����O3<Nv5�f,=>W��+I��gq)�$�@<4� ��pՎ� ^E���U�����2�b�A��砰(.�zr���q�u�,5$ GΫ��`�R���nSsoo!�l .� �$�7"�ƩRހ�W�sg;����1�S���#Ds�Ք���� 7���a_�X65 �LK���.&Osz��&X��'�h������� �ؤU ��a�6�MˠD#gf%[�a�f~���r��D���8m�������^Wy��ch���>ݚ"�Y�3\c
�~�ܻ�r#�M�.�y8�'V2��CC+F�D'�㠔+Ky���&���&�JMWIx��r�Si��+y/ g��.�C����NGhyK�+�ܚ��&��+t+��Ap��8[�a���,�~L�Z!�/V��8'�q���D�_E4��_0K�.LG��jy�b�/,C����/(�x�h�"Z���[�������/����g9Ӽ]r@�	�x����]��j�A�Q��;�:Q,��Lٗڷ0�!�a��$��[k,�J��>CM	@?���K�UL��mq�D��s��q� Zq�>�Cm�mv�����]n�<�҅��L����o�ot0��W�g�{`Z[^�n^��O����xJ���T����Eg�#چOϻ&/��޲���;(�B?�΅���(iT�|��*>��!���}�}�|�o[CB���y~�Ts6���t�չv ~y�硍�*!^��yL/��'I��叴�A��ʽ�o��Jz+��-Nn�4��t$T̆%{Ʃ��g���@A����b�8?M.�2�[�2�g�~yIu�!~/����u#SAR4����G��- X�l4*�S7mޅ�xD���{U�:���X�O��C�J�A�$~���'��T������t6M\02�sgp�����"|�J�W��KEV��qwHɪ#�6A������ׇ� $C�qN����R�p��"g
�f}��H�V�%����W#b�p�&RՊab�Cy���-J�=�l�aFUh�PуE����~�Ҋg��^|lDG&��#�p*I�k�x��v��׃�B��"�"��J���X�u�������qGtA(V�\�vكb�pv���h�V2�W�~�'[6�L��,=�Ȯό�Z�Cވ@'�t�w���"�Y���^��{����x�^<��f�}t�j; B=x>��T"��[�<��uա�#<��z�b�����)��9�:G$��,�
�ݠ���Xo��0o����>i�진�'*I��:�����2'�5<FKp:������k	�=�[`h���ӂ�?���,�.)2�e$
^�/��P�y��+mLT��>e�*���H�3��D�O$��n5d�l��5(��vp
T���Lgj��=��H���U�����<���h�Y���3�}1_��W��]Ŧk�*b)� ���g&���H�`�
wbeG��@K��[��������h���|�LՆp��j�Ѕ�BŲ�|(�L���Vz�~5�e�wA��@쿣2N��R�O4H�G�Pe��AT�+�Rw#=|5a�����^Tc5K�t7iPi��S�ߦ�4�Ȇ ��u�'��Xl�|���ۭtY!K�4��f��j7�0�2��
�P�}y�S*yvpr?�Z�����wG��B���=ğFtN]F�%��]�������8µ4\T[�@-���K�������@U/'��%3�I�Ұ�}��0� ��!��>�8Ta�]_��	�$n�����n"W"�G�H��@ҟ���Z)4-��Mj�b�1@�eiF}�\c\
 =M]����ݎ��h U|��H�݉�9*wh���WE�8 ���m~��������~-�`�����ОN��dw��8��1�Y���b�~J�jq��َ����ᡥ��e)�>F�^(�׹��9O.���):�P6c�'�V�1�z��4/�/ka ����Ҡ���ᦩ?�����<�kR0լ���6n���T�s��'��`d�[�'�(�+QDd`�΃y]/Z��"^=@����O�+�qr�8��� >�8V���%P�4w]/��|�	����QQؖY�0۱M�̒ S���nZ:�r�%�z��Y�"|q���vַ�w �0ch�AU$"�\������ս�� ���� �Xԓ�D��j'|�7gt��)�eh�x����2G`�JL�؏�`�L�K�@�>$�dz���H/;�ş3�U I\adù�3��͙�'��i��qjAg�p��{�i7�7.�k�Cz�fh��}�
���f���btTFpS�M�R*~�17����������Ƴ�wO�� g�'[��T
�F�%��� D�m����I��}����W�8�t�C�G;�9"�ł����\A�D�a�(=��sz�G�ԁ�g��]�e�b(t�nq8�Q#;�ۼ�����f�M� ��t�����v��o�;#�Z@�B�`�?,{Z4�	�5<��f�� ��r���3�D�r�M��:�@!��] uG�W���_���x��p�v��3����F��@l���_0f�̆�xV%C��dr�>=��H���'��'kY���}�M���La�=�3�E%���&dP��g��!u���T��gX��u~{C�]:0?&�[�M�i�B���5�j�"�R��]�MC���OH��L�4�����y�ͩ�?�@Ra���p���/�T*��( ?ji��5x{��)%��p��x�_��y�Gw_,������\H���_�~?�T)%���"X;�pi2��!�_H�̑Q6|y��	~�T�@'U���Vň
4N�>�V��>��u����1���MϬ�'`� �T�ן2�y�j��廀�zQjqF���\��r"'L��lJ�X��>a��n'�CU�u�hsq��3���m����Q\?b�Y<=]��V%\�}���WO�2dx�~��|N�:�ڧ���ExS`8�����E��Kq��L��"H4�	)�g��ݛ'�R���iŘ�q� ���ɕ��NE	��)X[�-Id��}��������h��)r�_V�I�:w�Hd���]�;��+݈��Wt
h�?�J���K:���,º�5�)��V�ѐ�G6���\��2�0�p�|�[�N ��Į�g��B��g޴��v�h�Ҹ�sW;SK�$yi����׬9��&�/j��W}�QĎ�p�r~t_A|X�/�?��
	����Lf���L��B��Ѳ{��h`/��cB�Jp/�(,-Xh)\7��Cti��zz��:k���<d�&9|�I�g�FmL+-uY8�L�&l���$��Tjt�^�zpH�)&<�=�kf"���.Ԯ��~���abN$ܰj�p
[��EpE.D^�I�/��^V�(�2N�9^�1�N�+-Ҝ�e�L����TUi�����F@VF1EO-{����f���Ex�<�>��F���S�#��oY�a��ݩz|T�H�T[��˫�N"r��gaڴ�#o2�N���+�p�9�栚��CNnl_)L09y'� eu�l����@8�VZ~k� =\�P�]��ڑrN���k��Ts�����6��K[��L=?.����Ϟ�D��dt�.��� ~ձ��+�QB�ԝY"l�g-}��g�P>�A�o������+�mS�&�M��N��*�%�$�ِ�����yv�Or�bƅ����
���K�����ѵ��e�6q%�^8��bJD�|x^V�cz��fbd�d�aY)�%�M(`O������H��N��3���u��n���/��:`_ѩ�����f3DR�ϣAb(��/�tD^�.��.rH�ux[ŮFh8dm���-�_���
�HB�V��X?�񾉃����}�+��F�m��@�˃)�+N9���\���q�"x������0�Ss�J��&5�P��*�z�!��+��J�AOr�Z��R `��|���%�<J�E.���>Fa���a���Ks�����H�%"�t�`���tS-�� ���\8�d���t(x�1���|��*�q��Y����) qD
J��6�L��>o��C`��kYg�v���o�,��"��� �V����q�;���N,WU 0ȼ��v�$�yJ�������Y�1څ{�gZ�����$Gp��G/@!�/�}��#ST��cO�(�̼x���?��U��aH��B��t��&�)
��wL�f��]BX*�l6ү�=p)�j�tE=B���u�����͌����`gzw$o��cR�2P��0��v�	�3 ,P8��[80�;���Eb��v�U���#�빕��Kaa���b�Q@~	Q	C�m�&ө(T��/u�t��z{]����ţ7�[�`)�N�$��9(���n��15���R?Ry#!���H�<7/�	o6ߛ��D�Ս2˶����
���[Gy}/�O�n}u����pK>�O����C�����RhG|��۫@�K���J�Eb�l�AGX*dfı�^�)����f=��@*�O��1�㌊�&]��2p�ݛ�R�݋>l��$8�I�~)ҫcA~TD3�fu	��;��b�4���s���*�X�4(O� ��8��v���;�}p��V����f�y��j���OSR�Yp���*6�j_�����=�]��X��ʽXٟ���z���}�WkV!d�{�3���@'������^�CВ1�	3*�b�%��h��	ֶ�.Z���7�:����q�o�"C\n�t4Ue2l�a�2\��t�ij�*Z�2���l��mP�����p�8X��'ur^���iL�����x̛v�MѮ����:3C$a޽̇|�d,�g�(����v�A�!�v}"�I��?���FH'��ͦ�&����TH�.�	j Ԏvl���5�(i��>NN�9���[�[��4w�f)H-G�L�s*���m�E�� (,$�Q��i��R0�㵫m�j<�6:��
�����2�&�#�q��6v��9�2�QU2T2 	�Lrq�!{���NP9�6�U��r�\�� ��� MM<��Sz1�/��VL�.-Z�:�����}�︟\�X�[VNv_}��E��V� ���k�̴z��#:����67�������G�i�������c`Ԗ��jC�X2
XlxV16EB    fa00    1130 o�\�����)M(U{r6B�?	�:3�G�wN�+��T 7��u�#��Z��;�y��q��ʡծ8k�����ʅ�i��9�b�u�.ZL �o� ���&~�s3���L��,�٦6���ü���0�A'|<�,�Y�g�e��5�1����Zc%�=R�Xc���~Y0,&����~�k�(�23j�w�[��B���E�����c�����=��<"^�o���I*�Za��x�W�����/�4�+�;�����ў���yL5�q7.��D^L}W;�(�φ�Z�m�ǭ�y�o�ޠ�F��(�r�w��z�]�e�Ȕ��q��	�Mމ��ʼ_)�����@�y�=͢\���%�(��M2�R�Q���0�$��.���}���T���y����5YM�S�(;5k�H���f��_K�E�I�<u�<*��'����ف5@�i�z�7S���J浅��qF������gG��7A�y(���erE���j�E�KĀ��ў��=�|�]ꦥAe�6H��������("��O`L�D,L�����n���0�ʥ�g�C� ��B΄�6��}�O��7R,���/�e{��c&����G��RΚVj�_� �FL������f�%�	f��>br�].�O�*�z�oc��E�t�������B�a~������DS�]V��)V��>X�I������n31,�!�JJބ��w���~nQ��4頣gn�Uu���=��mb�-)$�ύ�mPg�̚/G����K#
��Px��c��P��$�eh�WǿO��OBVx�. ����_a��Z�"|�^��9t�E|���M�Y V6<:}a�9����؈���O]}?����<E~�h����I��i��弳z���4��z��1���O_>O�
x��Ł-;@�<7�@�RN ����l}o3.(QD��%wت��2{�Vj�]߆e`�B���+&�!9�O㢺ױ1ԇ�"�FH�����-)t�����ޤE���$�`6�B�fX"�zK�ϭBWG�G�+0PPIR]�?�|�ꖓd��o�Y��SLB�@���x�1(�ֿ�h��H�����;��eǫj����Q�)2�j����p!�2h��ߥ���H��[h��Rg�%�G���������f���)�!
�w>aJ;�K����6np^��=�C����U���Ѽ}G�Z2�5�qԗ"���{���x���^&p��0��Wk�,��^ƪ{�zw�j�򵽠�/���A�V�+�-����7M��ǂg�R�� }��L�9S̃���v�%O�P�+�=t�7S��]�e8C�R'
0Q{�}D��Kg�C�pG��Խ��/�l��l�
��CM��N.��kY��*�J��,{���d�{q�����s��,�d�qD�N�8E��P�,S��W���m��o`t���Zf �%��Q�u�`R.�q���T��up۬��\�dw?�
� Q �� ��B��$@�Κ���)Sc)A	��oZG�����o+�����m�>��:�܁2c�Հڸ���뙼�d'�HRҗ���^�f���,_p��4�a�u=`g����|H��t9��ܤe���#�߮t�e	~�sN�mEW/b�Uڔ�s6�?��-�?F ��
���o.��oH����9c1�v����vbU'D�	�|���eb]�~�N�h�Z)�֙36�ҙPu.Na
�~���5qW,BW��^�7�d�⁑�p�KƘ���!����;�r}	�]=:W�r\
�� }�杶[���Of��@*�y��戂4�_lH�B�����8��.�eȄ�gM�z�c���"]@Kj3<�Xѱh=��?�<�>ˈ�w�<ə"���&��]�d�q<}�`3PY�'Aw�_�й~P��ߴ�%�Y�6:��nu�Mv��}X�g���=2/��-VBL+#�j�1*?�k�A���e2?5'�[D���LZ��\���{p�B�hv�Z���f���:�5�iQ�"���߁9�mӊ��RM���IE�Б0���s����|�D��tn�
��`��*�׈�B�uXR�s�힉K1廭5�L�mgb���|�-=G������Gj�G��ı{��;��.�����6c�MJS	�|PL��WV�nј�K����W]T&�%{�{�=fG��I���F��=��~I{C�|���(K8���ݛhcD5}GD���y��Zɀo��u�zn��3-�j�!,|�W=Z�{�~�9���|�X�y!@��^�M�h�E���ٵZ��a=W�����By�R�z��c�{��o��3i�r�\��]9?`z��,��^���S��mNhT~!_������lP��<�q��ɗX��=��!�H�y"����
��]bj0�ȸ>��)ZLU�w��W�VN���Z�U�`0�wE�1���=���������ȧ��Jw�9�L�:(���п�nv��H�.����t�	ƛ|��[Y+=�c����/��>{f�h�{:��t#�M�l/�*�9=h{ �n��[�� }P�F�=j�=\��� գ�<㢹�z3���7�TE�bpl_yx9]�����q�'ښ��ɢ���( ǻk�PʁD�>:
2Q������F!�xn|B�H��F�4� ���N�i�nE�j��@�P��|>�d'��ʹ�5m�Jo���ō�a-�!i75��Ek����w/q�T�؀�ƣN�ʪ0��Z��d���=����,��$�=y1+�G 	ү�������볳�\�b[V{�M�sʰH����s<	U�����Y�i�Mh��4�dơ�j]��*���T��G���W��	ݛ	��i��{��Hqa�G�`�����(�ԅ$h-��>��3���ۦ|�ݟ����?�*�ʉ:'�Kmʿ=�tO�yX�'�Nl�\o�2�DkX��^���hĘ"c������t����:���ot��A���ON��ŵ�`��������o��]��JsNI�/�3������o�+�7�/<��n\ģ���\�E�̀�d��$���~�|�pH/`��$R�9���N�0�'' ���jL}H��.��[���ffz0O!c:P�GV��Y(_ZL\���[b��;�� ��^V<�Ž����1�f�8��P�;�#mn���<?�aU-��H��>�r��e��'�؟L#v�':עm$H�|�n��dȿt��x;��O�HC���(�yJ�D��Ԇ���pظvU�T�}&�m�&��N���Z/*[K�O�u��&P1�lؕ@h�
�` ��s�v_ ��+j�1u�9��2��I���׺5�ꛂ�,#Ay-*��k擈Ұ���e2��V����]�
ҁ �Ł2���\c��?�*6��(o?��.H�ޯ�&+���FG\�F�VN�;�꩔�����܉�p;̤d�ۛ`cԸO
�d��D�|���Z����~ ����Cm�}���Y2Z�>�ی�����Ռ�E�"U�0@|��v	�O'֘G�����v���\E��/����F�WO������ �B�}�=̹��H����\���I���2$�&U����ftoeiI9�U��Cl��ܾq��(m�5���މ�Eԁ��aqz;v8?%H,�H�A_����a-��r��]��p"1�%�=��0�L&[��x$�w�O�#⚠*��S޳W9y�b(�����L���1��#���^H�$��$�4J�N���mD�@K������nao�h&����FG�DP�n��`���_�n�M�f��j�d��w >�ca@~��a�M	e����H��@+�����@8D,\@R�G9�z?/�eZ���D�tI>��A%Տ�Ɍ4����]dJ@����p�����[Z���m�{vD��Fw:b�c�"�<e7#���u��L�_�>� XU��n8���/v��m b1�vM�S�����~b���$��,W9�?�d���Y�j(����C�
�	��n܃ɿ�XѷqN^��G8޿�#�oV��ix>�Uk���Jh����7�?�����'@�Q���j��YP�?���T��D+v���`��b�4�o91<{�:����L]~� ���J������)����)�C1P��!�mfy�VwC��=�kH��c��.w_�>z�M"��ҍ�/u�Hm� �g8y���34�/�����<3J�:��w6���5�rB��(r6���+ڭOƜ���̺�z<5UJ$͉O�`����;�\|m^Ʉ���?k=VD|k�(_ɚ��;�r��mb��������	L�C<����x������H54N�XlxV16EB    fa00     e20\�/�E�g$sǻ?Z> D��z��|^��K�f[�F�{Y|9�4�<��<��^�S�O{0�K���� �K$�Q��D�َ�D׃Ȭ�ox��%<��2��_���c����aD�B��q��tgH��a��X��9��'V��(���'8��H�ӑض�{"c�\��s~7%ښC���2�K�tI3b�c�U�#�����:�o�G���oj��Az�"�޸F�u����w�[��=r�͹�����f%�M�g�ថ���3�mN�#�v�x�ں24�FVo�[B6�{?��'sF�$��wZ��^-�|ġ	0,����@�Sk��+V�J���m�A�{�y��AӢO���K�ǎc�5�m`!�㴅;���\{��@�Q�n����?#��`�Ӆ��v��=�I�}�N���6I����`|}��Z5�@��z���y�t}���P#ݜ1?$H�L\�#:^N�DH��܎��T�s+_]~�R�r����s��r34
��"��җPI��麸c� c�a���E1J�C�y���SdQ��e�S��M^��ćl*Դ�k� vi�|pȎ��uX�E���(1�(��6A����q<V.R���~\�T�Ƣ�������q��C~�h�������IrN8���d��5����4���V2�}PmV_�y���������UB�������ք-��Zdx��dV�>c&t�f���jK�()���C|\o���|YRA�j�^�C$��~�ԟS�J5�tƃ��Y��G�:P5������r�Oc��C��Pg�6�p葩�%�A#�	yIW����$
ni7�W��=�f�v��L5�RK�k�A���������^G���t��A����E �g��i%m��=�w��u���|���&V��	���i'w�M�C�&dV�ː	�V�l��m��΄�E�l�XJ�Ǖ�B�U��:������S��r�l�e�����r�֩�����/\�?B���m=~���OZ���/��С��bݼf�SZ�-vh�˜�g��j�R��N�[mаSby��;+�U�=��?�w/��/�!�?1�U/l�k��'ا�������ʜ�� -���UY]����M�y�����X_�s �aBhm�<�B�T�֞yu%bcB��t�������o����v��öp���3����(����M�4BI�T��K�Vc�pgʲt������P|����(��yJ�eT��	�-�)}���z��ѽgA�� �3�p�Kgq��PRa�đ���y�'B�jѽTO��I.F!�5�"�&٠ i�-Yi��8�T)AfR��v
�����c�z �7I��~S[?5\<�9sD!ifј������q0�f�K��)"�& �,���S*��:B�~u�[|@��������@�f�����'մ2wG�f�\��(�2���胓:�~�����	�P�Y��$X،�X�����F~�����MM}�am�}�f*� Yx�7�D+O���@�p���p�:d�%'��cB]�wR��c[� �z���¿�/��-7;s9+�0�;+/x���}�GfNKp�
���q`�4�Ilц=O��q�P�����G7��>hG&}Ì#D�
;�b-����A��v68E�Z�đH�a@�]�s�Y5v��ԏIx���w��0 1`�l����d�R���܃t
��8�b� �;Gi�^*DG)��������� *7"�����{�wwe]�ڟ�e���e���2�+|��6i2f��MF�Qܡ�+u�m������%�0��;��1N�U�ʄ�\��V`���M���D��l��|#����FT��_��d�_Ia��H����R�A�(행��r��rt6f��ǜXp��Hp0,%Ӎ�Y�PLk��1L��1�m�xޘ�Tu �̕T�dY�Z��š�4��|�x��U�(�C�@'��=µ�@J��7؝*V�a��g6n�֯�l��{�,.�',�p�G�D�
�A��"��u�%�T�$h'B��\u0sЋ���z�Ш��Bo���LM' �̸�c6����b��dh�Z�Q����.O���,45{�]	'��.���V���ߍ�ڞ�T?võ+���ο�f�y*��1��l�3�}��߻��S�q�gε����|X����ƠV��{��	�y]�����r�g"s�Ųe7L(Fs�av�:g�A,e.���͚y�'Q���*<�:u
��\���r��F��3H�	#ܗ��h��>~m�_?ɭ	*���=�ؽ��1�wU>:��MW��J���%���hKv�I�ѳ/�LC7�~B"=���M����$��9%�,s��u�Ϟ�ȕn��6x��(LgW44����	���F�!��_?���p5r�_%�e�C�̃������4.�L���!t���4ѡ��6}�E}��4�-�D����/k�x��Otl����� ��p�Ɉ._�sk��ޑmDu�	`k���wK������-W�05C���c�Q �7~�E�{��/;O�5$��S.G_�����,Ō�&��{�24��D���A�ҥ(����V�73�Hh#NL���cD��D�q�͂H:�ێ>�{Scz�d����.%p�@�R�y�)a	��_��U�_,qa��5>j����"�,k泟���	�L�?��pd���/��Yu*��
'"DI՟|�cVE@:M�?D�����>�`����ô��;�Z��_H��3j4rv�>KR|������P������=O�S�ti{�u.o�:eJ�[%����O I�<����j_����b��x�[��CܕY>^$ق	�b���%���<����}y�� �u��uZ�L���p5�Ԓ�|���ʸ�\�H�Z�� ��V�Rͯմ��f������!�e!_��"�.*D>��җ/����]S��G�뺉�u� �V/�j_̧�{.�����u���f��.6˽�ka;��qoK�{-C��^�d%�l�o��)�g^����B�lhK�[�F�Ru���>���n5�2Ij����ʮ��`2	ĪnL��l�p��̈ �6�=<�Ch��9;X�)�z(��x��y[b3�����_d��Ȩ�bRW1�c�߽��7����V���Sϔ�-���o�_�~��ss
zq?∖̥~����BS���d�7��o�Cb1�+��V�%��<�z��<���lD�Q;n"��D}`/Ap�{�SF��3�;jUNq�[th,���BV�B\V9ɬ�QŐ����kf0Ig�h٫��F$��r�0".����2$K�ZTb1�s)���g�|�u�C^�r,�(��ʌ���iH�cF�흧�%��&ȓ#������`�u���O�x���4�o�Z����3h���̔2�������^~��2��^|D%쑠�)n��#�S(BbI��d��a���n�˾�K�ա�����[�U^�RYPo��?,]�I����ߎ����J�T�QO]E��XlxV16EB    fa00     da0,E�,�x��G))̯Uq���p���غO��h,�n�;sD�؎U���K��1$���1���j������`��ю�A��E����r�J�Ff���8�v�x�����o��$GK�I���������H�a���R���,O�
��z���Kd���\`���&nB�R��������ϟ܉�(,��2��!΃�rN?�ַ&p�n؁W��ZQ�s���r��+�m���sH<B�0#�+��E��-�y��%3���X�˵�6L%�������q�b^��ji��ػj�ؕ����䈒����T����N�R||�{g�'o^���R��.�7;��?j#M'����[�e��Y G���r9��q����D��ˀ�!ʧ�j��H��{��Y|��t���DSE�;y�)�}�-4V R�6�����dp`�Բ��#�@O0�{2���2I�Vc.�d���I����rR���̭�����Qk�!:u��ߐ�K��;�s6���.��B�rm�ȧ����u/r,�*���4̔${>S�a�Y`�����"Qtd{�-��@~:�W�̚����M��r��'+�)@�xxז�l��U�TIS�;�(�ȬNG.F��{���N�w�v[���*ֿh�;dS#����:9��r{���sa�	���-�W u���?D�s���h� #�>�/��\�?���h%3r�x	1�6��T�~��t�%,���݈�rA��q;��X��F��f����iG��I2�a�-������f��z�c$e�<�i@�8�5 ��~��Qy�U���z����Щ�E���i_�V���g۲uC�pB�9����;�8���j�-���=��LBj�5����
��،	�ת�Qd>��Г�N~B�von�~�7��c��sٓl�u���B�b�vp���4 L}jh6�K�-bcs��,j�㻐\��:��=�8T�}�^�e��ƲF�.����]9/��R��U�t���F��0}t1ѝ��L�Sf��z��5���w�u�7��;�V0�Ϣka���$y�~�\!�r��{W���b�T��.�L}el��q��`3��v�����HKL���2��q� ��}Qn�OO5����[�^��՝��F�m�ߴ�l�DkV?ȢLhtu� �=�%����v�2ͷ5>�$j;%�G N�����p��Y|a2����>������3~}(ڳ\��QFH�10v,�j	�$L��� ��S%KA�2��$�2zL���Ӯ��c��ERl4F�p���vr����5���J�pvLED�O&IO����s�;�{�`�LXf��o^����{��A8��Q��?9UXۈ�8c]��,�1D�X��x״���l��wՏt��k�-[X1�	Tv N'ܨ;"<�%S�v�X�?[e�k��B�bb�]>�J|�$�.�q�W�78�\`��p�����*���/4gީS�v�`:�Q�6���WD�� �����c� ���I�էr�����T�O1�&b<ZFa�4�%̍`������k����n�|���]�&���߯�dU��}�\�su��<���,8��J����i+�6ob��'�Sޕ��]�n��i�Zɫm���9��gy�AL�0���c'�Bf�8k�� ò�&_�`C�8�n�����,�a��G?���,�@z�A�䶕 h3t�~��3�MϠ��DGf�ۂ
6s�"�"�2�&GX`ҝ�M��n��¢��H��Ț{��M9�3�uY�r��(Vd�,/<×e���om��=K������^�����LT��R��s�,6�">�)�|�^أ32K81��%_�$&�i�X�*e�Q>��_�v����3�w����=���xL�@���aK}���ڳ==��Pg �y��+�Jlw����qR��ںd�����S(�0���A7i��xsr����a�]Gx��G4cY�g�䢆R��W#��.��u��<��%-�?N��Uy�=n/qFb
H�gB'�%���Z���/]p/�$� uG� �w;�j���6�_�jy�9����q<�~X|�<w�J2|9fE>1D��g�d�wC��\7���Ce��A쮬|` �j-�ש�D����+��D��ӡw������D��1��+~�|-�����=�y���-��X��M�
0�\O7v@�ړ�y�����@Ud��w�W�q��M4��`�Q�������?���,\Vi�*Y���[B�o��e	_������7��ҝ�giXM�"�M�"��Z�n��(�ZS ���hi�7ù�iz� �v�P��I������G)o��PN��u�kA3��d�d�"r�Ε�tܿ�FNА#���P��-�y�+_X���l�y�M�FЪ�h�K8''�4$I�,�߆Me9*l,K�0�(�)K>��]H�΂��Mc)���@���AO�F�������M�b��<��S��Q����I5L�Phr=>w!_��=QQ=q��	GN���5��ɂ�x9Ođ,jd^���խ����-O0�C�L̡�ni�7�:n�K����u�>�Kq_��"h�>���4�l6}G�K#�:��E��N`�z�����L�Ť9�.q�P$>�6m���Ϸ�>0v6Em|�YC�����哣V����Q��F;�������%(i.��%\�%�-�n鉽�(��Pp�p�bi�&Q2�=��w�"�'���;�����!ܻ�,*�V��Pesz�@z��oD7=�����>��@�p��U�<�,��|r#�1$+�Z�F��u���vV�]B]P����0G
ځU	�.B���| �����!/�]��,'^�o	YH1�C�.(��E�A,�-�9�Nn_�o��x�`�i���H���&&�)���Xe�"ym��M�z,%d2�BB�����n�g,zrP�;.~P ن�]��i���u�f3����CN1و���|H+����|��3vU�ʯc��BЏ[�Ʃ+��+T�,H�]��O���c��NT��Zf�8cG��PuX�I�Z��ۓ���+gn�����rs\�pݛ��m�E��k�k�¦�w���z��_(R	w��M�. C֑�wr-��C6�Uyd�ߘk/��p^C�����^i!��St��B��eh�zYuƕ3S�"�L;s+I�vgb��ƃ�y�P�Rdi�l����;H?L�/�mh�l�h������OM��O��P��"����#�!vN�:�줚ݘ�\�(F�L��
K���mg�����~h(r9���ۡa�+�����5�7��uL&��Mk,^Ը�wv<���׭*�a$�]6�ٱ�n���Q�kn*;)������ڠHuHn�8M5��Y�#�Ia�޷�8�,c5�U/t�����<e�e���ms̾���W�%��\�	��XlxV16EB    fa00    13e0s_P���!06l1������M���kw�&��[%2sS��� Af�I3_Y����A�m��	&�r�7~ʊZ:���V����.ulF{��k�XQfK���䠙�Sc^s�h�O����!��D8����ED+�4��]!���d���4ΐ�q������[|@���{��-���;7�X����=8V��b�UyT�F��~��\�i(9!���Y��%(��-Lf9�������ǝ��Tfx  �<})�|ȡ��y���^��s�?od�c�$��b�Peiˤ�d�rC����T�-D����p*J�/�6�,����6���'������ezm���ɸ�{zk����!V�P���4�Ⱥ:���Qf}��{�s�e������6S0�>V�����2��^3�A|¥v��'_���
������_'B��d���o�����k����n�*J�C�JZ%�Q+�Kn��ǔ�	QRcVڢ�ܙ�;+6k�w���gbj�=f� y�%y`�����K_��Y�
꜅��4���p�,z@�8����G%j^hc��1����J�d������� �^BeH�O��=�#0�CV�B�W{�(L7��X��_%�'
 ;�/�7_>dܖ�:�*�L��&DZ������j��-V2N ����.�?�5DFrHsq��� /���tЍ�mޫ���� i����}�`I�����Z&[_���Ig��!���p�q��ڑ�=&��2��;5ɨ�3�bQ"g�K!�&m���vqV����0�lP�-�+�Y<��Cr���N��>�����y�'8�q˥����2�1yd�v��E��ᮖ��"٣�?sWv���a���l#[c�,���ʋk��`>-RR9��立�3��nKa���f�3�����7��`��e��]�up��'�V����]��4����q:�Ẍ́s}J�]�Ʃ��m��
/.���!U��e�[�Z?��. f���虷�K\[r̙0!�:3�(��J��G���w!���ً��Ɲ	*�J�SO1�P�N@��C����2~c��|í t�]~x+*

K�'-+�%��5��+/^��̈́�G-��ny'&�tC�(�K[|K�Tm�����%�w����j��n�oG{�q�jƦ��Xs�z�6ko�"У�c�XߌM���>��l�(��Vkg%c��'�w��5ornrY9i���y	���t,��p� �$y�o�B���䁛���8,|���҃ϻE�hG���l��Ͳ|Z<�8oJ&H�9<����!��@��}��E���R�Ârհ���a�}	�T�ʞ`!��Y'k"���G�����I�u��T��~�J�����S�,�>����g�V^���37�sh�"5��d�m�^XX�Rϕ�1����ȌNw|�0�%��X$��m��pgj�-�x��w��ƅ91!���B����.������.y��b����������h� �9�QE%�Qxg�X����<�d�T'�SFM�Vq�g�c���}���0H/�=9?�V
V� A]��,2M"�k�s+R!|QR�Ƴp%!1P	p3A���;/��\��#�Bg��+���{����e�[Ǭ�-0���ɲu7睲!�s�Ȓ��+[�Z�fc�k�i'�����aPxyH�+r!��ϜG���`�Q����~e�-��z��i5��q�f4�|\�T��Fx��#��&��	��\i��ҥɫ�\g�������^��˅*��F��"�E��@���v��d7iGB��n��=����Gn#���?�x��V��Av$��d9ˢ��O�!� 0�����}�x�E��j��[v_��X�ţ�ޑ�S�*�L���J2s-��$&�z�[��ǝu��ɏ�6����y�l�TI��+r��~RF�9v���l�2�躻�xB&&[b�K�ƬK�s���K�=�4G� ������o�c���F�z�!Bp���9Ncb�`y�[d���S�Z��g�+��o�@�͉��]q�r�u*&�B#'����tOI��Ϊ���W��N�Z��}���J�U��U�t��?�W�A�	�I)���Yď;�ڒ��#�qH9y��z(����tp.��=�ޫ��Jk�X@�n|�v���Ϋ��������"A���E?���~)}�u�	ܩC��"^�ǽ��;�Q��8ͺ��#��q��9˲F��4D�����y:�7y��B���@�DU (Ӭ���?Q"�A+`�V�M�,�KF��mDi�����?Q"�HJ
 [.\�
�R7��� T��;�qjz��񤊠���ٲ����� ����3ȁ�[�a,ԯ��℄�.����*���igi�:o־W�%s,��~��8��W��~ų�0ń����(a-d��N4��FW3���q��5L|���e�6~s��[���.E{ �	HH|i�x8U$�ܙ�[���M��t�$��Zeg���ϖO(t4��s�����Au�T��n�\�wW��:> �ql@��;������m��<_����'j�	(K��&�L���J=�F�h��Q�=`��1J�W�`��%3��XXqd
�{�މ~��iy��MY������s�� A�6v0��`�M�yiT����Cb9���=��&�ik�B[�5�|�4.
��/aA�,�i����p�)�ԗ���u�@�?�L��R]b<��������v�l�%Ѵ��A��(u2aYeE0���]h+; Ћ�+�̐�u9��+f����ޝ�]B'ߪ.�U{�:Wx���
XgL(��>F�
��I_s^�]<�^��nĺh�D��"@����1�?$�t�Q��S�
����G���7s��j�a����z������C��ǻ n�A]]��;tMh
�HJ�L=�%�]L;G6.?*ːٖ�Z��k"���P��;i]�ه����`+=���Ү�|��v-N �� �&��G�+D��̈́���'�?����ဍ��\����f�Hh�����������Xv��X���]�<��	 � �����4�%-%�嗡c���b�{�����^��
P�h┿�\�Πi~U$�����U<���_�a�i�ay]B�9�W>8�V[�����4�r��\b���y���2����p��5ݲ%�?s���� �~h�z�m��͏q*�l]�aZ_&�Gc��!q�MoӄD�2D�
Q�#_��T $�vl������Q��#�6���
�!�?�Wo�So����]��eZed��:���}�62���͡���8�\_cK �t"�V^هc�83I�
����5���6_��	v�ϔ���׽�v iRwSݴ�/���'Dxq������f%Bd���]$��' ��{�
u�+M0l,�ycwc�X~�at�oT��q�JAQ���JC�u����'�P�e��)W\����5Ƴ��Y��J@"��'Z=��d�~ Y��<X����kZ �'�>�A��UЉs�a!�!��:ծ���4.u�ո[�i(�)'TLGHw=�!�����gY�q/�F��5�A�x;s�2��c'k�r㖑eP�Rn����#p�Z]p����Æ�	��Ӹ��<���󊑢��6z�D����eA,'����j�bp�u͐y珿Ĵ�\����b�x$�&pL�m�����(I�ŴdZg���3�C��M:fq]��ђ�;}-5#:Ϸ�E�����L��Ȱ��j�6A�,s��Q���$�Xm���������2��7c�&���"k]!����Y�6Ng�G]zb@-m��ϰk�[�r�1۟{��C+���i*�J7M�@���]~�{A�|��;5���r_�y��Jd�S���;�S�����^L&Щ�.�ulE�מ��E�j�W�:	�L�*C\��tF�	��Wv�E��:]9��L��PH`�k���`l�0N<OR �޹�[5w�q� 	���v�ɩ�n��Or4Bc[��K�ǲ	s>(Y�G��� �l�ա���X��4a@������3+�K��/�;��g��Vк�$.x���t��)}u�s��7���k
���K,4 ۾_�aܮdܦ��%�/g�x�B��XD�M@�C��P/c"ITD?qP����S��8mr������s[
��V������bA2������ȣ!�B,54���	aC݊ 7���0�M������7l�f*"��+��R�VP����?�`�y�(zzs���~N��W8�K�:�H�[lbs�ʺ��i�)^6�+0���/�}f�ޣ��<��ډb�`�y�`���=\��d��Mۋ�m��TĆ����w��%����#ɮ�l�3�8��%Ï�י�P�
�PJZ�2Bvͬz�Vg޾�e��J��+�8����C����	�jB�����s��h0jI�$�E�ք�������i�S��S�:��W�˨[&
��N���b�N�Quq�-ƀw1���˱�3��˦�tdLCm,�s~0l5�����?	Q�n}�JK/�w(���ql�S%SM1���a�9r�\��ne�4=b�~��z�ڱ�0=+v)E���D��l
��:H~ʳ�F�(hr�Ǒ�u==Ac����,D��L ��K>��V����C��vzy}v���F=ܺ��b)߈��Dn)��n�����I����h� �L���a/@z	�¬0�6�tw�p�;"p#��� �B�U��������ٶ~��V��39�+q*T�1HG����<�IP.ݲ�.���WkN4�no��{��D��� �sJ#g�?;,�}ڮ�n��"�Dr�@�d���$�-­����g�M2X*��J�5�����b�>��!P׸=�˚�Ҕ
!�v����?,>.�B��n���G���22� ����A�R�љp�X���y�a�~��7����G��)}��'H���U�<0�& ���$mF��Y��o��h��)5����T:�0�!N#2��&���l�:\����heJH�XlxV16EB    fa00    1e80I��>;~~��(�
��V��s�}N�gm�g���w����Mj@�a�r EZ�"k吨��Z�7��vc��R6g��:冟�txp�	E���(�2��M�Žt<#��6J��o��M5�ꉼ?�Hx��b�%��qoA|>�)ę��I_t>0�bj?��h$�����μ �]�%&3�c\��]��*n�I�ܐ������ƕ���7�&�D�
<�ݎ>!<�e6�_�R�,q���3V�B	vT[�&�w��Q��)�f&mU#�?���.��E��SXM��G��Aqy��?�]W��ZG��Q��J���lk��Y�7�8*қW=��nh<�'��y�C(h��-k�e�v��i��*����7�W��b����d�7���7z%���_m�	�h�u\�3.��H?��UZ�z��
�*]�R�"�;s��=�K����=s���<!���[� s^c�s:�� ���M?���l��}7�=��=�U��_"�̼�0��rA���ӆ���Qt��;�4��-�u8C�k���Bd�
wS���o�)������I ��i�g�7�-��ȴ�F�t��XK��ޏN���^SV.T69c�_O��u�F�!f�R�L[T\:a/m	>�ϸ��CO�+���j����������D��Ӵ�)�A朅����Ζ8!#ʋ��� ���
�fo�G��=t�wP�Ҏ�B��Op�wNy�7
���v�^i_�Yh� >��Ckt�EAY��W��W���]n��la�6TJR��e�������
Q%e��FYͨ�xy��ڤ%9Z$�{����w���՚3����+�hE��Z���g�`��W4#������P��uH�bz�t���6�����@�]�M��kvXa�
y~3�U��"2���/1�V�t�`��E���/�d��G);���\���^?��I�Ř���Z'�-ݶM��ӊ��K~�A	��%���p�;�1(4/���̓����\�����59���bԛ�0��c���v�[Χ�Wk�sZ_�۴�qӕVRP�nρ5?,䧶�z�#�&�
h�����GvNL�#NM�kѥ$�W�f�5��^�aW�4��2l
�"�ݚ��|��~������rX�yza4�׌lN����KN�袨׎��%���Ts"���T��l��5�J��鼿��?�	�g~�l%���!T���f�MV+�|U$�`C�P�]G/Ghf�p�N��&�i�\߳	��1�+[��4y
ĦK$h��;*��sU�aj�ݓ�C@�%YZ�eE�=]%E$-]��Y�\r_Rj�J�s��P��j�v3�
D^N�r���0do��m�'�����%���5����������R��7�������%��B�'Ui��Bm��b0Xp��:�7Ɲ����݂k_��u��ƚ�]��ɞs��v��x�E���0���@*6f������D��������9T/:\��i�L h���;W�F9�?�{��O���:�6m$'MAŇP>ۘ��?�,�Tz�g��˝�H��+4�4� /'7���t:�P},�����'��`qo�Z��4m�׮��:0����SG��۩�T����/U*ms�㸑�R������8�4�FF�`�.���K�Tdv&��LZ���nU}�����RzlD��)��n��1X{LH�`
<�B�
�%ZQ�թ���Ex�3-��7wʸ�r=s���2M/��ս���b��F1[�5W�H]hy�����<�q��e*(�����>��j ��dV�����ש�qͩ��Z�������t8��@_h��d���%M��r���SO�4 G�UdJeƌLJ"�ŮUs`_{�0��zޭ�}�I�eM0�{a�A��xO�k)�\���$Y���03�az��璄��`E[b���;�p _ߨ����o����"���J�	^����h�����{�Ǣ��D�F� �3�vӨ c&�䳌�8���O�UI�::F�fЛ�V��e"���$�_�����_��Z2d/grXէ�����d��:��q����N.����I\mz8�����f_�&1l���xK�"�������X 4��t<���m�����(�2�{Ko�u�#[̈́��@��$�\� B;q���v�s����)�	58j�#r��BM��@,N���3�����Y�?�-�챟���>߃�-�`�թM��r�M �#T%���\��7��OJ�*��H�u�H�^�]2]2���iZ2��⼦'"y� �]j�À�b����p���ız�Մb�"�d,-�9b���!��4�^�[xGu�(���g�N�醔LO��-3���v��Z�r�!�@q����_����84�٧�'�9iTAlKq����3 ��W��WM�b5t��0e�CA���q�����U0��8v�h�m
�m�~Yb��W�͉T����		J��p�5˕j�E���Ѯ������i�Z������7�U~��BE��F p۴�B�9�4�� �qԲ��(�h��zj�SV�3�"n,ۛj��9{>k��\e�!���̳6��j J��K'��2W��'��;�7���$�&o�j���2c���9�:D��v6rW`����^C��o���f ���#�;�L��Q��m���7[��B@:���D"ׂ�_B	3��l�=q/��
dZ*⊼z+�V�i�e�߁o������(֞9X�q=m��� ���,���/�}~|�e�r���BcG��Ě8�Z5>�z�z]��y#8=L2�kb6��W�Kɻ�����pu�Ed���O��d����_-v&R�<͏8ٸ�����	�K�=v��r��O*��T���ce�A8��� >L���7��&5��B2L�K���C�0�H����*�"Y�"8�2��*c�69t������9'lY��.�/��5�FfqEq%f�+��� ֍6�&�������d)UW��'�1UE\�A��۴������X׽�h;l��Q@`l�稠�Y����\��`e�-D�x�Uj��i����CM�� ���|��i�[�o�4��To���;j��+��.�e����P4м`��3~�[\ˌ�x����a���Q�*�����v꼶�ft�~�ag$�,8p{�7�[�}|ɨl.܂
ѵ÷g98Y��q�҆S�!_?U�O�p�K3�i��o}�#����\A��8����.��[#�Q�UB�ua@a2�\0*�!m��ڝ3'0{�Q��)��|2j}�:Ӳ5$%��ckg9�X)47��5�|��=ʮ�����i�B�N*-�����$���Ē��R!V��L��k�������s�p0�k;p=ž�䬡��XZF5��|d�8\o�r%����+}���%��!��<�{���UFj���i�,T]^;ƺ��whu�9���b�C������\NS��B.�ͅ�!�*�ٟA��nB�T�3т8�C��̇�,���+�S�����C�C7@&�}$��0�Bp@��h��qP�#[���zY2�M�%ܭ��vɐ���}=����OZI���^4�Md{����(��"�#eC��&C�M�⤝��xu�1D���Wo�Mr�Hq�����3�v���L#N�!���ӾuR���d�g�w�h[��0N�ص�G�Jw��|"�l�Yi������AdeM���,
8��Hy���kz���K��m��w4	W���w�taD5�z�a:{����_9�L6&�X'r\��,DH���EI�R��L䖁����֕��.9yQ�?d.\��Q�6mo}R@w��`j[c���LU��m,�*��@�7��q�2m}��� �����d'�p�M��
��x��O�R4/u�^.���ٷr?J+/z����;W���zq��+	 ���E~up�����:��M��;D.0NI_�*s㟜xL]�hO��v��(E��x"��n��̌D;�IP������[]�����2�m_�Н��Q������O���/�&�����bõ��s^F%�C�߷�Ǧ]HZ�<��6�0F�8Ue10���Z�sï|�)��Odêj|A�P��pCT�mIl6롍f���#}��A�+�����(whW�����9��T�uh*5���kJm����<�9'g8dn�.}[���*(�M��&�N�w�jJ��&#_�҂�ⵇ��Fہc�����k�q(�� /v܍��FP��~��U�JH�de�G\H��iSJ#�>��pf4�K�Y��K~��π���^C͢�+v=	�������AIp��n�}M�~��|=_T�'��Sq���ܗw,3鎹"��ǆ���dfݿk����W4Tls>�{����Qh)ۀ�߂��n��*&	�GB��Q��`� ���Wݚ�a�Q71�Q�܈E+k%�'�m�}��s�R��ʌT�dWUwz�'S&�y�a��R*��:<h ��'[���b��
�x����p��Ή�kh��&�Â;F��g$�y�,�"�V&����o�`T?@�.P��gy:� ��߮����9�P\W�J����鱬3���uGʁ ��\�(m�P�]l��#��ͮ�h���,��17}���!/A��!����l�Q?�C�Z0`�ݎn䨨��N��w��fu�5(ݓ�s� �d��]�����$��"���h�����+�#�	P;~�;'�
�)$D�nU���K΋E�
򬽠c!���$3,w2��&�HUp�3� ꣀZ�Njz	>�}�'5��P�F��z��~n���Ə��:���Ǽ��f�D�MQ�+X�;�Hm�9�܂�_u�QW%PXW�ʵV���P�Bt3��y�p^��q��y���tǬ�%�?�f�7���^]��r����Q�t�tN� \��z��fB�[^v��5	Hrחl���B�m��|q�����	�:~:-+w2{������K7�\bhҥsE_&}:�&��OyHKl�\���*�#H�n�zl�4��ӌ�<<aB�Q,;5��m�S�JM����(-�������F�S���N2����6�b���x�H&�$T�ǉ�o���yJ���t��	��Uxݙ�������l!}� �Js^1F����Hr����[u�:C; W3��	�?ko�d�-���.g����*Q�o܆��$�(r�fʟf��n��`�����As}A���D60�/:��{��#Z������Hg���Ia�%;Ӝ7�č���tB�}��'�b.��p;�~������ARG"=�REt��Srr;��u���Uu����YTQ�f����z���w��	h&�c�b�˟�-ƪڿ�*�yѫ���C�&�~����Ay;���7�����{~�|?��w���`���Rn��Z8�XoAy�ʎ�>�0J	!��{����:�zp�c�^{`3��P6�^|EU[/nc�f���4��e4�Y�綿7�	�Z�Qkn�B�B_�n��x���~�%%��J�}�<�>V�E�QsE��*F��0Q��L�3tf�v
;���=��Ƙ�|C�EJ��*.[���R��1�o��]��	Y�^��gL��]�d��^����D�Zb����im����\��k��I�PJ��و�N�;$C��Z�E��8|��Oo
����ãfdˮ��bh�6],;�"=������4�C�p|"�� 
�)��{x�:�= ���9�C�l�P�=�u`W`gW>�4�(�P��k��4�d�q�Hd���ϗ=Ky�0��E#��n��sGsg���$ڀ#yO�?Z��ڵg�|��]Ú����[����]� ��5�[�zw,e6JN�$��k�zG��X�r�»F���"[�����ԫ�,(&�$�����t��Z!SPY=(�[Y�"�@�;?UK�ړT7/�����NI�n��'�7|�ϭ�o�� <U�9�Վ�	kz��\��$�BJ���(�+s��7Q��/^��{:([�9�:L'����/��C��E��l���h����kQ�	�A�I ��m�<��a�+�������j��_�c�K�,�V�yCx 	O��D�k�̫9IӎT��l��W��
�Op�hV��*4�򗆃ړ�[�ܷ~�SI6 Y<?uU.� t�5z�)W�.,:�)3L�%��DW,ͮ�I�\P���2=&�[[<��/=�<��s֖a
�O�ut�Ź�a�)s]'���iw�	�w�R� �@i�����lap�I)D�9̉� m^>��z�|�	���?�h���@ �'�c���q涌����:������%ǹ��0q�ZC_;{N�	���%��P�o	8U������d&Q���>�a:���&�3��&��S0,H�?sB&Ϊ�U O
�4N#fkp�OÉø�_�A_=�u{�LD��ox���nI{R�0݀�a*��z?�r���'���!��WA[����?��

��i�!���� r=�������<���Hp�pWߒ�֓�|�yJ���kO�����8J�������mr�0���ip�sO�Va�ϾB����0Djx7S��l*�F�B{+U( y.�=���W�狐)�(��������Pf������w�$�������ȼD����Z$F��M�GGxSܱ���O����>� ��q.������� �.L��Ӿ�� v]r �� f�6�u�w�&�k�����̺J�RC����B��mR֍9�q�?"��Xs3e�|}7�ft� )[�9��ˁ�O�%�Xo�|������п ��<ު�6�)Tӧ�}�%�eV���\���,@�]X�ms[��ZfA�Gvi��Nuw3�v: �9��Oϡ ž��j��eߏܗ��}P��CZf���a�����J��*F�;���7~��ݻOEǐ$�;(��˯;�ݥhW�v�m�4DO⸖Tێ�Z-	��$�u]�;
J6�eb-�'��e�#�d�d{	����8)��<���Aߎs���i�w�fj�9�6G� ߛp�cw(D3�稐D�mS;�N�6F��GrPC�h����Ŏ���Ș�M������[�S�D5��l�+v���F	L��$�WwGw�0[�n�� RЫDmo3�N���Y�1?BPV���*T�f�6�sg�t���}���$�v9:��b������=���7��?W;y�s{�����ǚ����tf��Ҽ��z��1{#9�̞��=�r^x!���p/t��y�n20]�{�s�d=l�IB���v����[\��be�@J����ix�,傝v�_��DE����Y��C:��u�ҩ���dG1L���6� [���-Z��!M��CN�̕s�
�=�dw�خ�7� g��_�� ���Bn|��y-jΐ��Q٭����}��>)j|/���V���7D�؜bd&z��b�%u#�����:w�n
$��ƯH�&��;��8�6��e��;��^m�*1"���cN�O�����ubm�tuR�{=�g"S�Vu�C�9NI-۲z\���Ե��`%��e)��@�M��R�8(-NmE��^`X��{ދd�0�;�o=+/��ku��.�5���Ɗ?��<��uHU�T��z;�L��H,;� �c`��tv�1����}u)'���\���G��M�28�L������`�k�����]��y�A�T#J�^��j�Z�o���H��H!%�XSC���YC�/*?�[�HyoXlxV16EB    fa00    1d20N0�����<
Ւ�i��KK�>�e�p/�e��w���'H?ǉ�B7�g���	�w�?�(/ఋ�d�k���|�J�8�茑���L��~���!��̉��K�3���Uk���.�,��N1I��y�ÞA���#�ЦW�(��d2�:���|��`�"�nk�ɒrț�5Q cs%�l^1�j��veQR���Q��c��J��.�	u�4���S��ƍ�:n{p)�-ʹuɵ*=;�lj}!�B���v�/Ta����y��҄ �"�5-Р�л��)J
�l,��!��M��ԯ�,��p-o���:��|gY�?4D}|�Z�5 �{gڰ�g����\L��V�y���F�,�$-ej�W�І�Y/ylo��u�S��������TT=`��P���<@PTy�`�Aj7Q=�1'A��`娾��NaCP"H��5�P1�I�$!�ݺ�@<ﴋ�ѝ�J�}�:f@�39B#�W}
� � >�!�+ɨw����'�r��>�4
��`���z��1�[j���A]��c�4"���?R�d1�h�N�ٮ����S��-?��y�>��f����z�f53� ����&�jMk��i�pL�اc�P�W��u���[��d�9�R��j��_�z���>���xe��q���	+Ơ��,�0�����߅6(��%^�.��OD������U���
Free��s�b��� wZWa�}@Eۦ����sʥ�x踪A���߳s�h`�S�#³� ��Ӳ��n$]R���ة��-Z�_��"Ld�#�L�+�@�^?�z��$4��ǒ�/�!F�p&�S�SdP"e�)g֩�pL��-�����]�g����6_8]�W�!�9��>��67ŉ��(ax|����|�:kI��8Հ��Kg���/L�_�k������TǛ�f�K3��!��g�z��}љCs�ş̦	y3����(Q��p��1ɔ�O���Ǡ�6�� ��iq?_O�+g������i'_����0�{-z:�]�j�H������c���P��|qQ����P_�Duz���)Q�I��t�:���z7�^eJ�c�~�~@�Ugl8�bp���w�<�����?��99��G�<�CЍ��|b��z,�hf*��<`�P�{���6���2��%>��[�R��Y'w���iEC�:G����U_�:�(�@�L�P�2뤶a �F���O[�3 4!��ʣ�>%e�k��b-�N~���qe�W�	- Ц���ϧ��S	��K.���:3�,e�36���o|��=�E��KP��9���U\z��"��*�'y��t�Q#G,i�on�FؒuP��s ,7jd)tl\�U�9�y�����B�v��b�4�9%�J�v�4�T�Iz�"b:�Q�+����k䳘?V"7	�R.��Kh�ӭWu�V�a�pUm.��͢z'����Ze%0�=�TKmG@f���1�D�?auOr�b�&�ɚ�V!Db�*Ŵ1jI��X��Ҥ�1���O>��T-�Ly�����	����
����uv�c�C�స��4��,�?�s����7K8�r�%:A.[���?�k1��l�ޑ�u9s�QM�B��'�놥�{��7��"��Y����c��H�1;8�����0�:���LS��3rw޲�$����zwv��򑾹G��1'-���
N�S5��L����V�1@��Ʉ���LF����u��<&�m�]���G��u"z�T�yAK��8�d�x�[����[f����O�DY4z,��d��7����6,H(8����5����	��|mo�ʪ��;�"����Z�5=i��:g��+9TZ���6ş�
���]�<��b���\�� �(5�ٞ۳5!�/��C[t���s���(�m {3@[��z9�$�zn��j����D��D�Z�]{�K'?��@��U��� S����G�h?0�o�*Yf"���I���m�-R_cdbt)QXk���<��t�  ���R�9<�`q�q~�������a'�CNd��y���WwpP�$��5�� ��L���ᙡ�,�G�i�D��������<�$�Z?���^�"��迹-&���f^Ξ�}���f Q�@�p-��L��PLr�l2҉DP��n�I��NqC"���ou��	r�/���>�#�
�Y-���������3�9�����?	",gQ
�����8\bnQ+Fd��!�to��x8i��)��$�$ 3�d�SoMA�G�M,��|ӳ����C&Qu��u:l+���"}Y]^R�a��W�0�?*J���hL�\�	+���Ip�?����DO�7�e4���X�4��#0P�[�:�U��~�ƓcȺ��<���|xGZ�,?z��@=�pե4�GO��6���e�l��e����G��R�P]�{Y���F��
�%gy�У��;1���_z�;Xp�S�(K�V��Ť���@�D����s�[�H��k��F-�ƅn�=A��B���]2��Lچݙ����h�6�Q7����&��g�%�n��]�����[U�qԟ����B�˲l��S�z�l`�s�_���@1��ֿ�4խ�YEָ�ы0m*�߱���t�iS���`��Q��cs���t"��������%���(�P;/mEXNؖW�u���l%���>�r ��8D
L��w��bJ�5W�w�lX�O��~S��s>����*i0I��TKs���k~�^���W�v�{���k� �O�D%�z�ᯗ�aR�Y�䃈g��Y]�]J>�	��U��V�/���Z.M��լ��9�B��g����������ӹD�@p.iw�`�b'wGphGDu�'�#��p�qj\!�P34�>�H9�-�]�����E��H�|�|,7%�;�:/����9r2�n�~�Y�E �d�|��jz�#��DK<o�d3z�m�rY� 4Od������8��<I����|��YE���0�`{��I���Ql��
�0��Ճ��-8E򼭭>d�[�ع��#-_����iC=P,���>mr�[�Gt�5y��m����m8����VaH��S�'4�F��=��މ�m�Y��|��Σ��zI٩���FJ�1.�!|-��_{Β�Erm�r�t!�=�H[�"���hs�ӑ=�� +�t�X���ӿ�1��ع��_8 ����#[�G�`��\�]�9��\�x��*jw \υ�ʚ~�<���~q=OZ���~�-�:u 3tf�r����:7�!U�=�M�[��=]dE���0Wvp���������������Q�%&�Q�X�X��p(m~Zi�F:_I�(!�i��j� ����#���s��M)������F�_��"k����N���@���e��!يS@P�qؔ�~Έ��%����+x���ݥ�,^�?�R4�}�IN7nnLºP�49_.6r9�.&R^�w�ּ�O��ָ�.��+�t g�4�#���S�)IQ�W.%�R0�����a��x�Z2���J��j�0�����KS�c�u\'���X��)|d�^6n�S�O�d�Vy<�����7��z����Ǽ����p���6�]8d�<5�̭����%��l=��5��\w�$�H
��ْ�:� �=�e��:���o0I���n�n��O�9�LI!���B�bXw�J�J�z��&6]���Vna�Q꽜�J�p:�����U�� ����Yg��ĵ��t�����T׈[Y[�	��rdc�����'�?葔��M4�F�˘f�w�6b��I��	D�)�(�ZR���Ն�-����o����=�AgR�9���x~�|T�l�)�%q���U���'��'o���Z@�,�Z��/Л�1��������������za柷���v�E�y}�l<���{RX"Lu�)dG��G��P.q�����'%d�RS��/E,m�H����c�j�y����)|�Q����.�{�Ѷ�8��z�BtG��`���j�Ed>�]#�#��]��z,g��k�"���=:k��đf�YQ̗_:Jd��Ntrc��٤O�6z[�����a�(�2	Vf���ƻ������� :�
��ͦC�@%$��a_�w�[��d����_إp)��Ah�����o�dD����$�]�6���LsR��ΪyM�¹H�,2�|Ě�,�^��96##?tS�_0�m���_��&�V2�"t��;D���S\|�;��E.N���p�D�W��3f�
7��0g��z�#�k3
� O�p�5�;��Ef�ðQL� ��|W�@u�Nn1��/��ћ�}|� 7}޲W"�78N`�
�];��*�Y�VT��~3U��Q��p|v�9�|���bp��q!����f���+��1z�jKI��J���8(J�x$�$�L�դp��	��qk�j4��q&�]���µz���1��%B�$�ߏ��@�����O��
V���y��=����=�_�'�|t�H(eo�Q	�K4!,?;���j=�V�}tAo��� tZ*�� �*��ɧ<e�RM��W*��X��A���g�l�Ϳ���I]*5�4�%r��aQKd�..y���Dځ%`w��4�� ��� �\1W��{l�*� [~_�{^+���o��2�d�e۷ƀR붑v�7�V�G�#@�z�
Q݆圦ve	K�C���d�g���ߞu�̾R�~�3��Xv���>i�?	��Z���-��ZR�b��������=*��аe�^����SVL�:_s�]#���n\�r�7- ӄ�c�u!�M��+�Y'#���VזfR'�`.��/<��<�HܷO����=����$��#(��Z_[�:�"���H�2��_IqJ��z.�=vL�$uT.���i�S��,{��&=�����Ԥ��νx�4V��8>r�O�:p�q4�7���y�v�O��'�x�W�~����m���!�'.i���BI;x�ƚ֫h@���7�'��-n�I�Una�I�.�IAf�<�b X- �3"��e�kwC���F��h�)�HR�B9	g��+�̅�a~���R�V?��G����H~���Qßx���.�o���K�zۡ��%�C(����Sc�͗!�$zbȸ��KD�B@��gR��x��5���A'������(\(�MU�F�k�y��??H��Z��P��u�MͶW�F`F���j얒6^�um��	�"�]���>=:���	�и#�TILB[:"��ت�bƍ�A��:?�5�HM0���ƪ�/�=�|�����xsU\���m3�{u�*8�Α6n�e$���b�AY���h�;��iG������V$�C��X�KB$�iӡK��=̨�nh�6r'x��&neY�:�\@3��T��w*J^��7�WD�`����I�iy6�ZA�J�1�����8^����O����SP�������Bu��D�F@`�Z-��G���V�@�!l�s��Ydz#��8�j0�4WXI�
/���KL��#�"!�\b�OK�|�����HЀ
��f��x��һ�c*�_�CXG�OdKG�J'��q��1fg�T@yF n<h��kA��(�a�L��":Zv�@��@ae��t�5�$��e��5b�->��U�vm��s��:q�1]�F�r������o���P��ا��T�g�-��
���^{�ldi�N� ��f�Ͳ�}d�I�������Zgz��$�#a��]��:O��"�B��7�­7?�&vC���y���~!��
M�ׯ�H���n���$6�Qܸ�Ճ��H9"����L;k�=�q��l�Eq'X��{���ј,(���U�kpb�}f/��t��vM/&Iu���n�%�S|~q�_� !T�:	��rnl��>�P��7hrW�Op�x�ۼ���͵���JT�xB�7�\�T�j�WvwKD���r���
��k$�����Ŏ���N��#�@�S�[��bn�V���/�_0Wڎ����_���r�ؽJh��ktBT�w�ĚP�*��V���L��Y{�#	�La�J��=���h��T���qhL��� @�e`3~y�y4��l�pѩW�A�ӊ�ν���Y��c*����Ş$V�`�[_���T��xm��i��}�F~>�
-)N�~�i96Qt�"[����U9	�����.o�ޛ�L��Nw��@���bI=������O�z�(�-u���t)F���W����L�=����Ī
F_��Z�@eq�ɇם0g��X��NhI��j|C9��8xۨ������@R��I>�x�9?����0�Q'�3 ��=�-8�\E���ګl���e"��xk�X�}���O��yp���Ԝ�d�/�;�ُh5�g�ڋ��֭�O��3�r�f�*�ԗ&[W���|�'s�T-S�r/�Yɟ
h�[C�T%ÿbe����_��^L�gic�u����'�gTr��
��(i,g���S�i�=8m�n�a�`X�8DC�¼��a��k^�қW��W9�� VWsǼ0֜堖��}�*2^ٚ�9r���^J�T�+
��Gz>��~|x��O��|=�S�m_�M5���YM�9Cz<�=P��9Ĝ��yE���hU|WHH�`��6�]D������t�-E�� s�oZޤ%N�|K-��,.5335F��j�.t�B,�R�~�l��?l?/K3NE�����OEV沏�Jopa&-h�Dۉ�B�/59@���/x�H�����R[$���S�mة�\m��q?_�K���3�ꆠ�=��wy�6t? $�%4�o�f����y�=�}F	�y��e�'�1�A�������2���.̪�����(��vU�B�~DXb���٣}b@� �I�D���&5D.z>Cu#��s�������*(,�k.f�w7����O�D�p�M��(�,T�d��ퟑ�m���K>k�T^���$�q�־"OHS�U��F����j2ҧ����vh�O�9�;��A��>���畒�X���-9G:$.T��n�tF�GZ�x�8�V�����e��#�6=���LdR�p6p�N���|���V��7p�qO��#��Qk��)��S�S��∸�+M���4逡�Y�ꢛ��3k7������זУ���]���5� ���͹�x�\Q��ņ?<ݱ��PV:~�r
��.�b�n�F�ٗ�{{�D̩%�y
����ԉ�D�y��l��E�V�����(�1�WF���7!?W�P����]ԭ��p���X�8]�hi�IK�Pt%?�p����Pi&�?��C�ְѧ�����UR��F�4�P�XlxV16EB    fa00    1670WiU��$`G�a\����~�'���Z��qVݭ	���.t��~�Y��A/���T��j���0��p1�n[�t[�����	a��Ly�)2x�KP
�Z���(��Ƥ�2������HG�j�H�X7g������W�;͞�F(� t����^���_V��I�/˜*��G�}���'�N�f���o�`�x�Cy&i��W-Zz��[����ic�[$q1��p�x6ک�џ�2�%+#ͼ�{o�r�y�ϿV�ڦZ�!���0Ie�\������`�>�7/w�M4���U;C�����o��N`�"Y��L�H�!{��\9ڮ��j��gl�m�����0w��NJ�ע���L�-ca��a��R�+��4�`W�j$�?�7�۰2�^&Sy�2��.�F5�x��DK���������$�~�1�:�yz,c/õ֢ysBxQ{�!������ yġ�9Ww��������Kr�ٳ��4YW���i	25�jEX��l9�Z�\2�g�,N��fi�����@��o��2@<��.����ƪ���#E@\^�
ω`+��K��i��Mt$��������U�+1ڛ`��H�i�S�~|�G���� T��$:P�f�?���#!7��4�=��)��Z���;`H�_煐9�c�_Ȃ� 7>And��5ǹ�X�3{��
�Q&�C	T�b�W�0�|�GV}0���d���c�&pZ9['��#�������*l'�ڎ;�C>B���61g(���\�e�(����O��8a��Բ@a~�dE���0_#���ӪG��l����ށ<���+��ЭD5�5u��m{K:�LOdI���A��һ�\��9Lz%������Q�RṮ�)t�<EA��@�����)yǢjQ���v0�>~{��
Kr��j���4�|�<���6ϳ'��Tv��gt\ĿkoEz�߮�l��!�g.��\��%��9��?KCrr�'��g� 苣���Q\_SD����KTTᯞ�=ߥ�Lm�82�{�l���FK��A���n��T�f�	l������ M��&;�X봩p؞s�}k��:(�7��n�w�
����@w z�x.&|��4� P޾�_I�q�+�4;ל�V]>��%Aʲ�I�c�eoq���tw�� �B���q�s��?�D���\E��i�����7d�2r=���#��)D�����2��.��KN�Ou��gP4��d�tw��XH�tR�^I^lX�q�t��L1�m�C���FH�wE�oiq�#���j�$ w�װ�ި%��ڏu����
Hx�0Ѝ�s��a�^AY �F�;�,j���^���%�{y�ZR�v@[�
�O[M��C����|/*:9��D�\����k^U��K��Ӻ$�Zz�3�����3O��19s�H��*���H<���$Ѡ�AOtF�<��0y���X��f�g�	�H*����2�(-i�3������&��*֡n�#P�����������`7+�c{�8�S�����ņ���ڱ���dx�љ���e=�Y�!��շS3%���������~���13&N��t9��e��Ȱ��OZ�H߳�:�W2�u��\�v{�Ƭ��2����4̇V�*�$3��3�����U~���q2��lٰ��w+V�Ɛ:��<_�N[���*yV��tUҡ�i�iAҤ�%I�8���K���zra�c�Tъ�s�<������t5������d�T���߿hVrA��jJ�\1��T���7���W�ؙh�[�ޮ&B�X���t"���o�>�m��<�U�b����k)Z����^��/�}<���1��=`
�t��z��� ���Wӫ��� Q���K�>D%%�Q�,��r��7#�R`$I9އ�@���1P5't֛��I/�]y6�c
/�j8��X���<T�C��]�����tK�0F����I(�BDް8��d	F����8(�`>���d��`�=��QB͑<H��[��s �!�j����������X�G�pɺa���M��DD��2�l҈��S�+r�@�$�	��8�gZx����i%p�]��4��zV��M��bǩ��]�yQ�+MQS�9�I"��K����Pw��+��7U��[,Jb32
��w���G��@g�g�X��%ɒ���E����2u�Xx�c$�$樢b�
��)V�R�<�ܓǦ�M=_�,e6�tn��QƏs������\,N���,��p�2`8���m.�B0A�T��!�5|d���ɞS^0���#��_�~z�ˊ���`��Hz�(��d�",؏�o��U?	O��6�����3F� �9s�Yu���>������n�P�^A�Y��]��!����Q�b]�#���(�J��)Yʂ��˱��K�$m�~b��[9��m���#�qކ�4��\X����s:����.|T�l�m�sxa�O���
{&��NzN���\�ي�����p "ε����>��Cym�a�zt�i�wa��G��A9�aN� ��T��(���_9#2^H߯��-f�"U��*q�	D������VͿ/QT����@g��o�� �v�g4��e�-�׊��8ک����,E��P�G.:tI�O�"���ͧM�g��A�H����2ƞ��Y��j�ڋ�"!>�_�6P�nhT��|;�\j@�L�)���ݸ�̉[�Ѧ_�hJ�(�~�-�L�D��ֈC��g���L'��NZ !�&���DMkD�`_�8Y2�����|����B/M��c�������:�@�PU~�eL�����0�&�e��FH�^��$�+댰�X�A���c�M���!��0w����w�ޔ,�{ ��&���p未�z�D��q�<�}���bS�Rn���"B5�2`�Hx>L�q�D�{��Z�fE�b��k�C��؄[p�|���Fl+v �g`k��P�h��t��^4��@���������3����3���h���HBgіe~�}Nx�@8��������>�:{��Yr:w�b'���l�c����w�C��!SsjƮ���,�r��)�3!0U�D�Ma��e�W����C��:Y�}Up�Z��_�lM�Qa�Ö����X�r�o�3k����(��� �F���VG�O����ZΖ��D?v���<��i��7S�'^���E)M7n×��3�,�NP�&
Ty���-r���r$�=b�l�}��;"������ϢM�UL�Ii
�9�	�8cd�M�~ŏ����ͻ.��*貉��F�2�5�[I�bW �CZ�����0&�"�����X���e6���߃_�ZA��H�N�%���]'k���-[���ΐ}q1�fȞ��X�-~5�
n� %3�U}oʀ��&����o��u5�#�%z���5>�ؼl��,��Wy��~�G�gDb	YEi �2��/?@���ˣ��o]��`4�uD�Q��s�e�9�.�}�P Ĺ�6����L�4�P/����Q���I㊣�K/���M��o��R-�����
<�աrdg;�[���fv�~�``���a��� �*��������H�}c�^����0}��k�`傑��ީ��H�)Y�C�9��]pկ�,6Eq�C8���u� S�z��Ĕ	@c�E�@e�Kč��+�)�Aj��SM�eh���\���4'����T�%�_�.�#3����⊾���u8��^n�*�V�X8fiȋ��m�C�?eJv�`�.�:��C��1���S���� �z�w1q��AiE��4Tv�ތzz<�q��_��b��drZ��I��F�>Y�F��g,D�\���D�*�h?�%��W���O���=��W�6�H���ת>JW7u��xd\��<
��c�1]q��>�=�$�T��J��D�8*�Y�ڽ���ʃK?.��E�1iެ'�vA됣?0��S��>Ys$��Ց��q�.�ZZA�^�N�+���9�	o�.���нx�7�1:e�=O�(Ga��A�Leh������R SE�]~$#�!��e�W��"���0�l��2Bڛy;h�/�ݨ��ݐP4ѥ�TA�������`1D���e��鵐�E՚Z#��q���
���e�t�h�Y�Q�H��9oŚPF�_�BL\�lE5C[6н[%Fzu�coi�̽s&�z�x@V�~�vc�芵���C+S�EXM\ Z�s�Q\4��r�Љ�W�d���\�.�M��`v�NᚭiU�+��֨�&����/gj�Դ�<�}���c������?��p g;�Bݾ��ǩ���A{�w������	t[�O��a��������?d�w�(�7�����I4���[����r]8�R2<�7�R����"��ӔxE�i��H�]4`v�����:	�� �M�VB���ڌ�9Ќ���Pe���G� \q��JĂiS)Gym9��\����_�{q�^Ba�e�d߽��5]ZU)��	v��14W,[S������q�E�a5�-�G!M���7[�y��i(i�&>��/s��z�'Ȱ	���D�J���	�OO1�I�8�#v|�{oG�,�Kqyfr6(J�/3����qO�=���$�s�wSV��a� �+��C�ay�,bb/3-�GG����)��]��qp�E����A+���E�[�X+�e;����@�F��[���>��=�Mn�F^r#�o3Ɲ���OO��y�<� 6~:T�6iR��O�m�؝�fQ�E�ت��HA*Vۖ�O�^�l��fHp��R�H�	�����S���,��t(����02%���P� ).�J�տ�X��y9'��πL�Z��RdL̅�Ϊ�?��Г�b�	:���I���m�����
�v�$7�\�#�O��/Z�٩�R�_9<	��=W�З��k�r�T*ѣ���J�E��ǔH�'�CY���a�W���v��.�~�� q��uMEW�E���O��5���7�r-;X�k>6|�b1t7HQ"�3�zR��-�"�PYAP6�Gԥ�U�$U��U���[M���/#��1��z�)�ұ�K?��D���n}l����`!����[a	;�d���{��zi������Y�m��U��0j��d���&׶W�ؒ��Z��/�}рa�F��'qE4I~�>��	�i]+Y��-��c�j�>�oU�׉e#�0&�-zڀ�Q�����1���AQ�Wf��ûӽ�p#=�0�T�о�n�w�LA6g��|4'�E�_�J0!a��>��h^��4�G/����론���L���!��#� z
t��<~8��CF�,��Xi�jg3�UӊQ̾$b�@����v����K��� �<�`�����_'D��L�U��YzD� z�S/>�m�JB���R�;���庶��O0�G���%�=�\���
��d��A�V"\��Ldu�oTOM?!u�bo=Ũn0�xg�:�0:<�O`Y`�[�I�-37v)�
6b۹�l��4�!pG��JٻJ"*��9o�s���o�W���۞1ϰ���T_�<�)�� ����.~��6�M�O��/KN�[O���a؉�4B17���˙W�H!Pf�
���#¥XlxV16EB    fa00    1740Y�]-G�]��x�a��Y��������8��9�+�����Gt�@��^�c��om�.��w��\�T����Э<JQ(���uDK�QJ3f�\C����LAK���D��@N4Q�k�ϳm�E:B����,�>j:P�>�*��MYh�
f\uB�T���:�G��~�*�)aD���o�pz n����0r���S�HS�Q���<���rS��`����Fq��W�shymgI�Vz�����^ogZc�is'&e�Iz���
֩������6A9�W~��2��#A��� �P\��?|���˥e��D:��Ы[�>�p��و��{;�ٿ�R���s�f(�%Z+���H��Ƈ�����B�0�MI�诃ml8�|*��G_W�[v!�E����lҏ����A�y2¦�ګWM�_�sNgJ�*�_�����98ʤ_t���=I�p){^"8�{�485�?�@�?չ�4�L����k� ���e�
�=�@�.6(�ޛ����#?�x�O�ѣ�5�\�gJW8���Yep�B����f}߉Q]@E�9�"���j�I�ۿ��6�����@Bڱ�\�ȵ��?0�(�x���=0�����bhgʡ��������laކ��v�z@�+D����yn�0Eq��i�1'�`b�:�=���u�v22��j=U�Cg#l�?O����1�Ŋ:UH;ί�0�W3��P�T��C�UXL�B�.�T%���>uq��g-��|�;�u�q_�u�Ľ���`VzЩ��&��^���0c�4p���z��o����"�m-�.�нN+�g|�D3��ŷ�V���� ��C Ɛ6�#�1Z�O�c�q��t	l[ԩ�q{
B�R~!������@gt���Э��d��� ��e�������L�/�1K��Jt��!)L!f��ۍ��A���G���P$X�Gڿ�AU)5a`v٘U�s��a���	��o��A��T����SZ���- "`͞vxˡ����HK�u��k
���y�^3?���ѝk��m���D�f��JϏ7���+/_��SP�N)����0�i����ٳ�)#�acӚ��F<ˊI]���ѯW��$^����jW���t�p���^Z1�sh�����X6,�RZ=�Hb���&�	���M�:}8 ����@6]�v[�8滥Ѕ/���	�����8B���c'�P���O>�g�3+��m^B%s�2���#�Bܒ��?���]���t��V3f�٦(3y|�?��Z����Un����ĊW.��=-�����w����^:�����7��XB�o�����?�, XuG �HJ����9����V�N'�yWj�e�Z���"��aK�K[SÎ^̸4i�:� ��$v���G����-+aHIrWWz�P#e�t5#�䚆�2OG�[�;��NS_A'˛Z��rAH��W�$�<������w�@4~���A��0�2ӻz;�� �B�R�Sl8��|#3�a���G�PX�䑣m������_ɯ��mV��vV�Fu'�ί�ȹ��0-������@�9��-(���ͬ6z�E���R��҂T(X��E G��h��sX�_VN�j�%�'	�����)�Ǒ����49u�õ'����w����dPK�B6Jr�xJM��Wmlcjl�v'5��
��gx.몬�Jԅ8��K>�1D�~�*�I��4Ն�/�ER����o��D��&g�%����y&���0���f�a_�9��CJ�X����|{g62̣/����n�W���q$�{�v��7?��
�h�0���/�/6~�f^c�.���_��!�DY��Et�vY(4��������'/�-�*r��JW�M�����ɜ����77B%:�1�`�ʖ�>�AoL��s�I8זn�?(&�~ʻ�9��M��J�������^�5|�W��{��ݡ�?䕕�������wR�F����W�<�M��1��p��,D��v+D�|2W�*�)�3�!�]����a�����>g�Zfe�����|�����\�]���ʫt�(�۪zq�@2wƄU�V��wT#Ow��]��X�����/Ի���}Z�B|�x�Y�mn�R)�p���N�K��[�؜�[М¥�p�&=8�o���F�":N���d���|��!^Q�<�Ҿ��Z�z�+om��r�[](�U&4�)�Zp$�H����;�x}�m}�1�WrWI�79Y/�x	l��kd��Zz�'�D�Q��\�5JT_>�� �9��b��N����A�]@� /{�f�5�VM ���E�ü���Ѱ
X+aX���I7���ç�[9PtN��/�8��W��'g��,�s�������b��~�8�������P�>_�g���d6)���{�Y9Q��^��?د!
�b)Ex�g
�]�f����'p�u&)q��o*3X��`�C�f}o5�m��ʃ�'��?�R�>�ͧ��ڤ�M���Ŀ�CAt~���� �t�
���k���3��g�NR��4�H�7�C>�!a��vo����b�6�ݵH������ N.��!�5,o|\4��߁|N���|%$�l�:��S\&¿� cf*;�8�,�0��5w³�]�h&K	ޑhd�;č�S�H�p���z��;���G�9���: O�i1�Gs�8q�X̝܌_�Pė#l%�Lf�7Q��Hf�Z�M�^��������z��,�=�V��e�?��Áad�Ф�E�_�K��d|�,wn���-�����W�{?�c�b?24%Q{�wh}��&�M��bCd��b�s99aR��9����UM~�#*��ʱ����E��7�zr*�B�ǫ} >6@�����h�'�%�˚S�85P�F�9u��� -z{V��,g�t?S��ޏ_3�	W�5ϒ��=G#v�
PxL��g�70s`L,@���)�����<�f�I�'%����0�3������~���()�0}e��)���9-|D�`��w�=Rí��g╓��	1�a}�C��4��奣4�>ly��4	���\��t����\&sܼH��*���� �ȈA��^ ߮�qң����PXW�h���9ԕpv3H��A�.�ߛ$ڍ)�{ֆ*96�?+L��j��n���=����X�[�`���Ay�_	R������=!X�G|E	A`3�����.�/�Xv������#�A�'E�r�{���QV*"Xk5�&���MT�$�<�Q�,S�-XE������5ؿ�dv@�h�3��c�0v�p�Z*�`o�e�"��[t��C�N����}ĺ���N�/���ܳH���R��� �|#h��I�ލTMI�#�_�����d4���v�i	cuQ�]WUP{?p����v�SVv�~/+��&�@g��[8e�c��c��w�Lb��Z�F����!R�9\_mp�t�q'�D]yq�i��!��q�~�@؜��&��[j�Rr#J*t-��P��cnu�.��>EgQ`�=�
0�� �}���Eq@�U��@�l�j]."H�*�BPI�`�2vN�eƯ��*�Ca��?��L\�Z6�rD^�>|�.!@������g�߮[�(ݗ|���s̖��=o��t�KR�rhD#��g Դ5�d �6��֜d7�/�e��`���[��q�̘ꭤ�Oj�<�-�kq�h�/ER�2�K�f���b�Bi�#�G�ńM�gM��Uw�O�m�NħE�5�<�\y�
������լ�*:�L�ţA�.�:N?�����[g;���Zi�*�����)���\Q����=�E�$�����n����gS�Y�С���^�I؛r�1m*ˏqn���l���V׷� �Ô)��w�rB�,6�)B%��AZ��_P����S!�13 ��;���m}����k���6`uԎSC�FA�8��c���l{Y��UU���'�fI��'�!w���f�~q4Q���G�3�h����a	w���rO�UG�G�a"�=��<�	V�u��0p5��x�. �nM!x^H�c#��z��������q��ТW��Kɺ8�!�����L�Y�fp��k�p���{��Ͽ���d5��V��K�x��Wh���]Q�#�qk&�gH�9Mw�7ӥC&��K�4ۥ� ��&a�/��h��b��P���9 %~��_�Z*�F��P�m�DN�B����EEɰ�	�4�g��5�uZ��0��J�?��u��ܝr[�e��Wҧ�;��n4�%I�kO�&*!��z�n&��#�!��L���o�	�z!ہ�RR4�j�0:����g��:���ICʺ?p��4 �ӓQ��#���`�W�J��s�tw��Y���3�$���üp	}W����)�
�h{�
g�G�����$-�vQ�d��ṸQ\tif��*4g�M�DA��:�������LՅ�]۲��uN�$�FT�`5��D6Nv<(�r�un��[�X�����O�M�Τ��C�Z9�Hr pJ	q��:�8�ʐ�Hb7�o��Iň�!�,�.~�b��p�b�m&�~`Y���,�J�����T�h�3�
W�ٙ2~�)��|H�*c�3E*+4�PGL\l�W�����V:��Na4Z5��+=t�b�^,\����?=�[��o`&#��'=�E���~;{��UF���-5d�4��]LE�(הּؾ���(��ȯ�i��»��ׄq{Fg�jG��{�]D��teT�n�s-�|�<u�e���ᚷ�ګ���ۆ���C��*�a�bp����ǿ��&Ǌ�~.y�����2��j��7W�$;��b�b� \ }���X�E�>oK F�[c�{��[Aq<�W'�݅x�3�X�e���-HDr��Xs(5���AzQ$�4EA�����m��l)ib��2�Y�Z�b�kP�#Y�@�ꌷ�F���S����8��lJ*!�%��o
i	�v�?����!#BV�4�A����E���Ai4DC;Z���Z�7��Ь��b���-i�^�1bI���)�P�Ӯ�P��m��l��ї���j�zB��G�'��V��5{)�0x�0��&q��ug���\��*K��_,i��M�-�KsǷ����}�ϴ��7�e6J��C��^�Σ�<؅ds�!�uЭN��(B�Xѓ��}����]�M�a���A� ,t�٭����Y5ѭr'؊K��A��Z��J	�ԀDKk!������Kq�hT�S��^֜�-�ԂC��~��ӊs��1t,����F� �i5�K.���l�#W[?���ϼ;%gV/7�i=l�!���_��x�Ոʐ
�=�k� ����0���|���ˎ}�pA�p�g8-KDwꪝ�a,1�z���������:`��I�D��{���'�z_.���1,S�+�V��#��欺�I��'�h�Qv����fI/#~C��$zJyO�)<��²A�r|j��-�g���A����td~K{�}��5�v�3�G<c�2'��T�ޚ6��S�Æ�vD�a��K�����l�A�Ж��kC���, ��B��5[ā�t������#�-�o�:!a��L���w����	�4��7�`݂X��ģ�Zk� G�C�t�E�auc=��Z�����X]`�����O�e'w�����!Z�Di;��W)�X�Z۔iN�&Eg&�\E�����l�>���^�珣\\�q��Y�~�3��':�L�^ݠ���r, P�\Kt��o��a�4�:�=Ǜw��8�[�f���b:�}��g��/��
�N6D:d��MN���h_ܷ��vP�2��^�r��j���*G��DoXlxV16EB    fa00    1380l�s�ǉ_�g<���'8�7i%X�F�э]`��;�v�z�N�î�[�^�����l�z\!#��vً�~���i��T6�@ӏ�oDD`h@�g`��&ꘂ�"����ߊ��xq���n<|_߭(�;W
�1^ř�[Uv���l�!���Cz �n��J5���@}�5�32����Tb�>�2[� ;
4��x�g���ރ#�ڽ{?'Π���8�0�Y4��%ĕP�f 8�Y��g>�6�.�	~��6����1+6�R���g6�k�Ե��)Q��Ի����I5�3��������x��}"l�l�p\�Ϩ�kt�JT��K�X����w[�{䧣h����"�V|�I���Y�:�#�g���k-��ف����[��g:�݌��;�����y)a�N(?����hQc�y_�A��J}��ܰ�NЭܻƃ� PT�M�3��Ӯ������q���H�j��`�"3)����Z߬���ݖ,.}Y[���q�t�� d<��l/?k����f��o!��h��L�톱�=(�խ��6K�K@�w��R��#����s�R;*7?��S*��� �sAe:���iP��m��t�_�i�~t9�P�rz+��8���M�q?Vzs\��3U�t�J�)��V
a{�o���?��E���z� 2'��"�B��������3���	�p�.�j�7��|b����j>�O�N�b�����ZU�;�y�p��UC�{����㫄[��q�����_�_Q����آ���2�dW���Zٕ���7c�Lww���"��h�ې�1
@�6�7��:�Ӓ�iJ|]	��z&�Tn!�`Z��F�3^�ٚ @�j
~ތ8n��.�Wf��'/`H�!j��7T�c�N�	�{G�W��S? ��r1Q����8��,�u�}�p�����#+r�7��獃�'����-�bF�(���պw��gCz3*���}�m���b����Cx���6�eлiq�e��<�"7,�p����#� gH:��1����i��Va��s���F�:�//o�o+ld�t�t3�$;�,ų�kw�c�0a�r��E��� $�H�W.�o�E6n|b���`���(���?��_"�M7e�c�c]��V3�	�r�[��q����)V�q/R(	�)�)"��H=�����|΅��+�h�o��kEs���Ek�7�Y�����p.�|G`��w����c9|���:&y��s�����Q����{�&Vמ������l�&$F�G�Oe�����^��oN$7>.m��f	��rkgC�,�#��t8A&�p�k��p�/�9Da�e�ʠ���TY_��o�?���� ��{�ΡY��R�s�AWՖ�����\�XI�3��a�r�F�Ic0�����1D���d���KG�>�E�k
��r*�	v��nRݻv]!�]��a���-�w.����z�~��V�y+�F\��w���`#�D����R��C��B�ox5r&��-!J!Gi�׌U��d����Q�U
��?�C��v��z�cx�	�?�e�'�.��C�H��>��ħU��b��Ge���"3 ���(��$+2o��)#���-%�\-R�$@ei�:�1"����.#`�\��E��HK
;tō{^��Ҏ�7|_@�d�g��֬�p}�nlL6�`�ih�����f�fŤ0�J`�c`ٔ�� �T���N9J7�M����$�maf��9�k��3��|�`
.�Е[�^� ����'�ni��%�"�L�zp$*i;i���y�v#=D�)-\~(an��_�'���x���ϕBlÂ�G��~�����{�����Y���3�'���t���@3O���aT�h|^�
��c�8mS�=��G����'"��P��ʮެe����a��3�<BG�y�d�+�0���.�x���N_���k�Ε���TJ������h�����>�֖of�M~g����)�Q�GP2F�\b��ۈ҃>W��L��>Z������y�jd��8�ܩ�)=�I ��50S�/#e_�q)z�{Ԟ��F䇮�r4�w�[<���k-�+����~����{=
6�d���<y#�f&�0"��7G׮�29� x�<FW3&��gVSw���)���V;6�Z���q�K�$Rq�ܣ��pt+W�V��F����}�������Z�p�.�\e8X�d��8>�n��K��Q�5�����X�n
�ٸp�|G9�H�p�og�q������{������I+6C8h��	y���������]4:�P�x���tîm�J'=Y��q2�(V�
�L&9{��F�_r�ee�~W���B	��0V�{<YP!2�ܼ����2�K�c�h$�/�w�:b+N�4z?ުQ�cr�[�̗�'��y��Q���S��R0�E��{:r�+5��I���
�x@�����=����.N�*�!2���9����"�L�*����n��^�gY�ְ�u�H��������ȅ��~���&�T��k�aVU��<bpM� 0"�c@S$l���+ۤG
�:2�d��!$V;���#�${�	���cN\yqnta+|��1н�>��1��cy�B�'w� Z�5�Q�&����^��C̧���;���m=��;q���b���2��r�{y4�F@ yɥ�81��f-��&��G�p�X�
Ϗ\��D�UΠWKn3t:w��}z=�z�FoM$ L�'z�D)�F��z�ɨ�Y�ROX�%�d�rj�v������� �^Y�ؤ#%��DJ
r���6UAt�����!����a?�R���ld=w��7TE�r�у옝�HRu��{ �2/�)�ݐ�I�\g��K��((\����G���m�7���`��d���6)M�����9���t��K0#�ݴ>�:)gX�b:�~_K�*|�p�捹ʒ�?�Q�(�����q���<��|�&�ع�jh�7y�@�g���U�f�,:�[�Q�.A��s��� ���pb\5�����*x7�+�5�O� �k,}s~�i�N~�U3��%�1��8��������A	pF�?���E��W�Jc[{K��uV¸V��?[e�����hJ!`J(��9k;}��w��Q7V8�����2���LM�"�M"�o�.?�G`7��w��׸Jt���M��k@��Q���H?s[}*�a���3´nOM��C�ƒv�zBǸ:���[�Ld�{`8��O����R6���y9��p��˒&J���S��m����������	�7����J�{z� %s�)rz�BZ�r��ۉiq�v���G �J :���~�f'�L�W
� <� Ӑq~߫E�qi����SYeI�w巭��w5qR���R���1E]������\���>���kQ�d`/ڵYaz�*]��8�{��r��v����u��XG�lP���L l
w���:�<:��ut�U�tI����W�6CD�M��D�Ց��&뜀�O�hЊ�d(�ք��-0c� �t
N忦��M�U����D�� D��{:XG|fS^��]8�7�J�U�zO'�Q��<%����W���g�p�~�A3)�c۲vQ A	�d`�K�r�c�9����	&�a�s;C��q��2*88='z	�S"D���"+�@�KyCC	9 3E���i�AŌ���G��I-A�C_�I�Ά�������9�'D,k8Z�X3Xu�y��ˋlr�1�7(�Þ��,�Q�X#��~
����W���(uy1�kCʽ�]�7�-�|g�z�r��#��9����j]΀�-�4܀�Oa�J�&F��[���u��0(��E{�H�g����$�m�Y���g*�_nq��(���M�3��O97�I�h;׊�tG0*pt
�MCn�G��2�p�d�2v���Ƥ�@�<Ƃ�-�8��킦%|��J�H^N��)-�8��Ӟ�Z4˻�y�;�vF>��G��b5eu��j8��A'&Rm�{���!@l��3|3��p��t�/;�7�}�鴊b���B��W3�rX5PE����a
�ܟ�VF���B��4Z�����lD\x�d�7um
�'I�l��R!e#���J5���A\��Q��^���V3���?	c��xϤ���y���݇�*�ht�K��3VT��\�٭�ߞ̑$���h�}�f��Q�"Ύ�f8��s����8/t����J�ה��b�S�	��cܸ�MT>.����.<��s�&�C̍,u��ߺ{v� g����x���sEL�����u1X�Xvc0��Ԩ�x<�;����x��vk�R���2�0�Q#$��[��s�Ҟ��Z!��(��_+olz
����	Jk�&��eKtl��孹=�wDdEZ� �G�ȱ^�c];����/)��3.zm�P�n�f]���(G�g֫R�j��"Ծ=16e�D'z�HE�B�l������z��K���A�ac�>��~��H�z3��t��s��$�TC�8	~�g%=��"�o#�lM^ʼ}_*��=;�[��	j��*�>W�%�r�i��K���%��u�E�V �*l[�0��>������-C���wwDT��rH�^�H"-M"r�Uz|�J��L��pe�l'#'2������+�)��V8����K��N|�ύ�Mʸ�T�=v',�û�Τ�v�)0a-�6<��|���4�s^3��g�
qI�u����c�4{*/Z�Xn-�H����z�3:"O%�<�F��)�U��`��o����ݪ��0�8�r��R�g��J�}�G�F��E���%�~?�E�J ����!C���Nn���=��y|Rx0P�����f���+�$�s!P!@�K����j6 �4j���N�9�|v�XlxV16EB    fa00     720�2��V�C^�Jd��̿�o��{rRw�M*�>+�9��'J�A�{��CAC��Ц Ӹ��# �	tG�}���9\�N��.��CjX�`韾�W�8W��B�[�9���[S0pvy�[��8s�*Q���P|f��3�U�ݛ����#Z�1[B}g�`�)��(�n�ɬ�i�,~�Vlվ��yR	f|�f�W�Ws��3=q+�Ay��7p��Ov�|���&��;����x��J`��F�+�gZ�N�%��PB�"��^�:��ȇ٪MF[ku��������&5&����L���/0&8i!���	��9ƀ�Lb�A5C���;���ɲ'��z]�ňR��!$�{�����R�3��&�t�G���rp�y��/ט�=/�����nGQ3?j���(�g�>��ʝ�	����#[�J�\� ���j�e/��;3�ϓ��j�r�.<��?5IX�8ϒ��F|���h5���A|�үc���S0V HK��h�
�94qe����2��:�7Kp7`��l�A��GJ��8�RL�g�����.�-�)��ɒ�Ka�a[1��[J<:S��c��ٳ{��K�O�`�T�`]��ӯ�X�:��J�K��M�q�aXC$�9$�����h�S��餸Jٲ�?Bh� r@?�� �&��E��7Ͼ�u�
��؁�|l�ӕ:�~5�K1M�H�8�*Ud�sAʰ���S��]J��9��ڥ�`&�.>^�:7|�D�c��i{�)K各yZ�Q~���i���R�^hi|��Kov��G��i$�$9��T�<`�G��{M�0O݋(�yˊ�>�v�ɭ����x��dQ��������C����
C�yK��3�BC�AoBF^4D,/���P-�N��G��rJY1��R#h�\:�ݞ�s�T�D�lBtcݝ!*6�Nh�!��{y<�ϔ�炜)8n�R�I}nT���3�D�N��"�����rA/Rѓ��x�7��R�,S6����zo���o�t�<�1Q�~&�����6��k�߰�yp�#}ǢK7}[!�!��/����s�R�P/Р���ZłԬ/��o��7O�G/�h�n��N|��O:Q��2��!^��Q��
^�F�C��$��I<��L�A�:-h5�"v[�����>dH�@��A;\�?W�x0�ݑ��ᠹArc{44���z?>��:��⦮�~���	;W��tC`Vs��;��m��?�<������u׮2d�?�����関)�J0~���0`o'�ߔ{LrO�� �e�ϟH6��!���P�RH�_v("K��ٚ�#t���OQ_:))��5��v��bp]D¢,k��ii�Ҵ���}0��-'4RŬ��I�YMJ)?�R���6���8n�����4�P�v;M���3u��!ߋ��)�Y�QFL�f��00�-mY�q_j�\�)]p)"=��7�OK�+y���o�v#����á�_�m�*n�ٞ�%O�WN�i��DP��PP�������Hxzx�m� v|�Xb����ȍxQ��d��ŐfIC��e�ъ��q�{���w)d�w�>��|�c
� �C�$O�l�S�7Np�oP��L�P�A�d��`^�4�E�2����K���oF]�S�W����:���3�7�q��'�GVײvd�T�ȹ_	�B{.;T��[����0a�NC[���Z�,�45�dR��	>�j+�I/�l�K{ZH���gXĬ����,P�j"���K�_d`�U�ߊ�`���$z��!KnM.\RT�~ʃej���[k2�:�>V�� ��[XlxV16EB    fa00     670����]��FL��w�^�m��i�>���y����J����A���Ϗ��Ӓ)w�������弿q��C[&)�H�|�z� ��CF����@�( ��ɒ�U}f����_�γ02HhE���͍�"S �q�Dx�)j�&`V�Q�B�7l���-����³`�47�U9f$̎���;~9��ܺ*��5��������	"�Mpo߲�t\ݨrRJݡhS_S�+W�uc���S��i��k��[��ظ�h��"�t)�,a$���F����@�°� +5���	h4��gҢ�]@
k�Wr�n.c�g��p��xӆ�"�'�1�t�/�0�@�b3��<S��=nhU)���B+���g����g��̛e�$������������wO�����t$"���2��,��s��Yuú�"���d�='V���E���l�/�w ��7��iT�9���@�}N��Qx��I��3�
=E������+׫�s�ԍ:]!wA^���2}�sبwG��JQt;w�8�@�1	ű=��\��)�O� MV����1Rܹ_��TP������KTI�A���L��_���5��>�9b�[�r��]��Lc����$�a�;_J�f��C�ô%jzٖ�#�n�2!�KWΊ��'j����#ɕ������e�"�����7Hj7���E�#��)GQӛ:�����y�lA�m��Hь�R�2��|Ep�zX� ��)�O��?p�������׾���]r���|��H��� �Fa��ޠ3������/(�p��7�7�m����x#�u�Q�@i��Ɇ$_���y�P�,���q�D���V\u�X,)��,��ny�T��
QC?�PG���6vj���Cj l�@��'|�A;��T���%�PJ�ޠ�A������f<���.�������\,�kf�;�+Y��VY��1�4��V������=���q�b��������R=�:c^��^��BYC��a/3�$܁��G��T��;5
�?�-7L�����'_���2�&�%�Ɩ(���3��6�~�2bs��� Q��c�:Ǌݨ7�9�E���������#%&u��4rG>���8�~As�[ǘ�A��^I�%툈�m�O��[1�@�3_��=�*��J���ǂ��Ҩ��]��}%����b�8�����P��ɍ7p�%o!�W7IE�P�x�*b-7�]��]�i-`!8�i!����g�<�"����k�5dv�`[�0vs]�Q��e��s��7�v�s��M<j���(�;�K8yG��>դ�p C��XSߙ�UFD WV�c���?����$V9vE�Y�R�}#�0I��A�ˡ-��k�+�\��Wy����
�q�a���/Da���n�*�Ԕڿ52R����$L�j	����1x�s��"^d�.z�2�������E"�}�!�fwQ���m�֮�C��6n��ȶ�J'N�� @��h�;_ꞁ��CU��(���'`n~�x�:G3லTF|������$�]�42��;�	9��I���k�F@W!�p"�f��G	�)�� �(��m2Ѯ�ZCU��Dp����Nq�H�!'6��Fgզ��[�碕K�U�@<��XlxV16EB    fa00     590��h-��ͳ@a�}����n�_����)@
W=��m��l\{��8I�Fn�[�;�����kR�ă����,ލ��n���y��K���(�z��B�wDćqq�X�-5LoZ<��3p�>���k�Ea/Cr�&�Iױ+�6��>�{N=K�<�xg�}̆P?��m!0����.(2�L��p�XZLʴ @y��&�K�I�j]ƿz� _�f�"���ླ�!q¹�ҍj��aQhi��(������zKt�o����Hyr@�gG���2ި_`xu܈n$�Z�X:h�vklKa$FJ���r��-V�OĴŔPeGK�����G��
C0�	#nfc���2U�m�o�œ/��q��/�B=�<p@i���N{��ъ@��p
���=�7=Q����K�e���v)@;w���������T6�,Jo"�ӻq�z%i9��Ӂü�Em���Wt~ᓆo媣��T���.���7G�<�6%��iw2k�������nrp�M0����U�x���z�.U�m���Ƹ2�z	dȂ�ڠ�-�ў;�bg�jt�lļ~��?X芨,��;!U����{�A��Uu�u�|')}4�a�*��8J�L�~B�.�ۅ1EO��G�?�X�WA���|��!���VeM&�Y��5��(x�������l��^Α�>��V�[	����@m�<��[��*"��ský?壗�-�<��Z�~1%>�� .5��q2�{t����Z 6ڄl���
 Iհ1��t��&����U��og�,;e�� �gGf�/`�X��5�p�H� 6B8S�ʘ5ԩ"7�����5�i�}��4�X�� ���I_�.����6�L�D������1���!��?����_�
L̄��E��d\���4x���P���dl���%�j�ŀ���xV�biWn�z���`vy��Ҫ_�*�_LF��%j�k��أ}3��"͈�<XqH�tj081e�
J'�U�Q�����˫�x� w�e�m���S�ǂ�F;��0w�$��'-c[`��웼6�,�܋�G�p���n���N��߃@�@�O��Y�p�$�@65������ʟ��v3[��76�DFO��é��}7Sڏ'��\�6�y�ͮ�]�p�Rު<ܖ\>S��G��WlϺ!��D���t��h�m��Z�Tyh伙�n�r�纙�(����<�c .�Flޜ�)k�=f�D5/� ��Tm�P��'��S+'���-�;�`��4�R�Iڰ4��t�����5t�yU��@6�+H=;��^�S b�`��'�"���!��qE������'��ID��Z�.����tg=�&�1��}��3�Q����e��&�x��yN�*1Si�v�C�[��9yؽ_v�Sm�Ǐ�T�W�����XlxV16EB    fa00     600Jm�^1����,��]8r��W&(���cU��e��>$��uB�T����S؝���^�@�K��U,��5�飉o���R���;ԁ�Y�ˁAc3#5���3Ao���v�:`��%�D���	��{m3��xV԰�Fr���� �X�
%�b��&�X~�%�h�d����S�����4�׾Ϩ����ځQ�O�����>C�}��[q�G��IKj�eEy�iS���=��b/��&:N�КR
���<�L.U�?iZer��6�l�վ��0Ķ�	���L�/5�Rvqy�x$iSf�ʓTT��pB8ֳ�Ũ���{;��CBM�����|'}N�񢇌���(F����9-�����c>�	�����&�C�l��[nTv��ۧ�H�
���u|�t���5�.(w-FS=�J��n�yhW_r�t@"��"T^�~gM��� �+9��-�� �l	PY��EYaʼ
��%z��Q �'aga�UD� ���3A�-@;o������d1�QF?h��;?��T@x6g[� [���-Xߴ]'��l���y�^��y��˩�K$�U�@��@���]��Uh�T8(�����1����� :N�F��F,@M�3�W���[(䊁2'��V[�!巳��=&2�n����#�]�$���,�s�~�Y���(��q�#\,��;�VH��^�x\�!]���FsS�FY��烂Y㏟>���ZI:�67"��Ze	2��|/֯��E�a���ί�6��ӗ�ju�dk��R��yx5�$`����O�?���1 9fEz'�t˹�;Z.E�Š����&օj�	Y���H\��u��<F�R�^J�Q#*ؖ������#��4�����g�׌g(}E-���^�x�?��8V��f9!�W8��?�9G��)�o��_AJ/Ϭ���Fwz�d���lM��b�%4^nXBc���qM�����
�r����P�l�b-������#.���$�Z�;����+��g��Nlb�����4DDw�)���Aja7g��{m�VCl�kzp
��
��#ڨ#�jm��j��1�1�YG�W�o�|AZu3w�^=cו�|Fj@�I�WQ[�C�P6
�p�|]�<:�cSj�$���.12�<g��Q������E�{�r���opR��Nޟ�<H������#yYdH�
�+�q+c�Ko�"�n.j�R�q��
��;*�=�/�[%授��w��K���%�mRd=�����������_���jQ�lҒт
����f���6�Q��N��$;x;��%a�#�{-9%"~��`V�F�NO�"�A��y��e�Ł�ře<���$���`j�J����^�fn��"�<fΠ���n�g���<���*Lc	��w,��s��Y�䛘��Q���&W��r�Ѥ=|�z��Wa|;�$��u�8��o%+K�[����/�[}kzr��yK�B��*�I��y�5�]9%ǁ�=x�|�"��!tcte�Y&ʙ�#�0O�25�XlxV16EB    fa00     910�C�r����(;Y��_���9�8�1���}��%Zx���N!�v��5�sZ��-H�Ѳ&`Mr`��c��U�k+�����f��q��B���h)4�b؅���<{�8\�kj�ȡ��n��#�9�M�G�3������־�L���{_7�ɚ��֩�Wi�D��9_����E���J

%"�.������NK�('<�1����_��uo$Hs f�gf6����x�X�v�Y��q�AĢFQ}3�	�Z��1Y��	�h������{d�٤�X�J�����(^Z���C���y3�霍�aW�s�OC���Cs'��z�s7ճ~�X��Aj�*�Ƨ�䬙�,�V}�v^駓��|Eݬ���k6We�۫uc$�2V,dv�3�{���Z_쌳�������Ԡ���ZGռ����#L���#"��+��if�;�F���$ጴ�Q�Y#dҩ�v���� L��J�093Y�Y�P�R�,���J@�GBbN�[�����H��b��9_��0h-?���'X:�u�X%7�e��:��3�~���P^�1��g�%I#,��w���,��l�=K!�*������=_L�R�
�Kt�?zFj����{(R���z��o7ǘ�"��0v�aD����ɶ�K'j�U�3�ͪ�^���g6O�p�+ݥC0�!Db�0lX��'��:��a��T�Bo7�cI�� � �u�\�C�vܣ䀀����H��_�!m{��h�E����v�Ra�����H�(L�OX�����Gk��{XW��)6��{m�k�'kΠ���2�}���/�ef� �GX~:|K�7@Kk"�eW�c���n�S��� !ź�y�;�~�?V�?j��2���� 쉚��p��]�w�0��)�p���Pզ��wu�eq=q�7[,� 7��܀ޕ�Rw,'"���=�9*km
|�}�\��D�D=����4�I&�M�r���~$�HB8m]7p3!��f��]��
>̲�yg�~Aؘ���$�f��7	�( �L���~w�	�U�āa�����J����A�(����P?b���Z��7��%��\qWl�^�r�7<�
(��K��$�<������>?'1h�k��J1
��s�z��c�����t���CM�(fb�Z�\r@	�{�W5��$���u�6�ZƔړ��hAɴ�*��V`����i�Z�Ra��N��.0�w
���=�"	��9V���%��G�2�+���ޡ:=x3�;�t�@�&�%�/����4�9h���Q���n�^W��s�+/����WÕ��K�x&�dE>N���U�6��[������D�累A���2C{�4�`r��� �)���&�o��R,�P�b�jYx��cj���=>m����$~�ͽeY5�#�A����ま��A��k��������4�^�!�M]��B�����4���a��}���=���yI$JYzH��-��~%�{\��6�$N��&QR�[l�h�j�]c�Mӈ4�Pֈ���i�-�%^Z���@/��V>K�����(���ϨQ���EͩG,�Z�Z��P�R��+�7���}C�I|_%�,�G�J#��|\ku�w#d{����
�sG�BmSqE_E���V��T�b;ޟ�z�![&nh��xlJ��x���0g�5�hM �������N�-��z���5&(�w^4m,�� �/�"TS�G:�%k�"�dE?':Z:�L��Mip�R:�e�%U5�p]�aM�J�I��Dt�ڣ� V
�}��2�շ�\�9M�O)�H�u�b]�+�18%T�]�~�Z��6����g	�g}g�;5��ʙ���� }�4��� f�)x� 9�L�<K��H����ech��G�-��ٝukr��j�sk���r76�\,?o�8���",�T���)Am}��cE�y0+��\�n���
dl|CP�9sS��E"�ul�	�2w,���s�DȚ������E�S�u�b]�9����r]~�����9�:l^���#.cCd����[ ��w�n�v�H��_-�v	S�@*����q^��N9������(��;��:t�(��+oӼĠ?�k
7�S��e�X�T�&#��n��g�0��0̉?%�V�7�JRtRR�)�c�l.��#.��v6C~ߏ�PxTU�W�b��2�L���]����~�^��X�0XGt�Fu�v%h�۳����y�ୋ�;)8�3��QQ|���"XT.�j��L?v���O~��x�A)al���d�UL��#��	�D^�!*t]�Q����t�s>�7�XlxV16EB    fa00     a30@]���	� e����S,���"���-�IS�M���B:���VY��m5�����&sL.y]�^����e 2NMo�
D��/@�cv�IJ$'e��v�Ɲ�dx�g�,dΞ���ÿ&q �b5�������'�ň����@L��K?�yL�U�%�M�L�ʤ��w��m�MJ��}�3�v,6�	��1v��2@�>��0�f9���c�I{�T9	A���}[S��4"��Y"C����4�19�c�7����G�iW.�DUG%�GrhD[灭���]۪acz5�-1,T|���Y[V����'@�Kp��-Dr�!�@��ֶB���(T���,�L���d�Bo�����HTϟ A���. �{PJ���p׭���KF�Q~�z��r�?aE�B��s07�+e��wL�Ml�j�oާ��#�K�d����7���8=P�� �r���3"w�	kI~:�i��ό�aY����ۼ+m�����M !cp%t�(aC=8
W����]U�fM[uz�� :�{Xq^3�q��-3k(�A¦ʣ�`�<��)z��ب��k��[F�䛾�M-�+��V�i3�3N��;�3̇�'ԙ�"�K�4�[V�a���sTS�O @֐���z����"|�\�~�x�(�v��;��J���Z��u�X�D�W��`�%�ϒ��|�s�ấ9����oV7�x��Y��6��g��<-o1�@@T@YEe����2| ��:��������v\m���bl\*r�:lj��υdև�B�8?|�Y'��L����|�O����wypT��vtV[�+I��"�<?�紾?4�X.5��)����*Mb���i�5|�Ύqw�Z?�)#�V�.�-Y(pb�B�S@�1c}��7�.h1�9��6o+7Q+:���Z��h�-�s���V�`5'�J�ᮀ���W��;������{��K���Fy)��@6��!��`я:,-��%��"-\���ʮ�u3D~,�|IX�����U���.��(��_�/&#v�ޓ[J	�y���9}�LN<{BH��/�-�<꧙�P�(�+����W��|��A�{��$H�^;[� V�7���"��k�l�\MQ��<N6�x�Mc�:�?�.!_^M���ٓ;����c��M�e� �̟��؇w`I��0��`�rf�n�)G@6������'�t.�=?���.apDUg����,�W��xYZ��n�R8	��u���G�^X��򰗓j�MC��2
Aw��M���G7�uM�t���*B�A��, E������^��Do�O���<�؄<��b����iJ8sl�1�Eb#�֙��H��6��9��^�e[�@�}���2�h�8A�P�����;,��@q�-�4��Dwx���р: Kl�2�c����1��ʚLb6Ry�ة��a(h����6W��3y���/�[��� �{;?��6�v���/�"�b�S�1I������<��W��s
�:h�)&�1*웰BfI��G�����劯<'�t,��*���D�;�҃s���.�X�����a��'�y(J+%	6&SzrW'Xs����pt$�<6Q�/��63����30��}Z��d�����IT����O_bG��UƮ�~��|�W�`5�u�O ʕz����lw'�iXX�;9���B��Z����gFR�y	U !��j'Uo(����~������~r�4�B���׸��`������
��#x	�X��WC�5��R�>	�I��+���������&��J�	��M����%��n��q�)��Ƭ{�D���Ƞ��)To��l���K�1 �3�v�_Rs)�N�$�H&��#6ɸ
�\i�k�[V�K��*����,�J�)E*T����c�.�!�!<5�l��7�/�\�ɦ�|iC�3���1a�2NO�ꗫ)F�����P�����W��/8��Z��p�sWc���L���RGY!g=��PhR9�f���E.8p�OĿت[��k̶��y�ȋ�y[�G���p.覯Ҟ2��v,\��e�����gz��PV�{�$O�O_[�:�����>��"��e�T`X��_o�ԁ�Y��,!	��P �[�-X#���p4�SP�&���b��У�����`L�Z~'1�3�_3(x<VC�V�K5)�wc؍a�G�|W���H}DuN�빜+�$� ��2���A7��d���"���'	i��ʍ�ٗ�!��,�4�~�:�0�?Y����Y�FvA����8L���1�
Ks�L~�
���|�N�=s�ʍ빖���^�e1�����3dzeG���i*g�u�]
��6 5�Y�:sQ&f�@�gK�S/��[q�� 3�ӱ|���������Pc��
�5?��0�6�h��/��|/_i���W�=u�U�$>i���-���|.�H��c�\d��Κ_b��"q
���*V�wҠ�#�LfU=��N7��h�"$��~�0��o�����ei2O��	ak��D���H�9�s��g�J�H=��� o��oz����CԈ̆�C�s$?K�:���(XlxV16EB    fa00    14a0\�5�5�2�Z�q\Zγ�_�2X�;�"2�,;l�C�}$�#�O�W%��R=��A�Xsq�:�0N�=���Pw��n�"��|��ɥ����_���}0ˋ,5i�`����F>��|
��)H��KZA�Q�a)����3���R=�Q*t��vB\Y^�v��Д;��@/<�/�)����������7}+p�Y���T���+Le��~\��
�Y��H<Y��9�m��,[��aY�0��>sw�x��0)���T����8h|���]�W)��cR���c���<��2��Ju۠��7���=2��%��&*�mq�n6����Jc�"]#�뙙a�Uwv�.b� l>�`xݑ�|'��ސ�w�<�l%����l��0<��� Έܖ�
Y���y2fm��1�&���s|Y��o�a����q�֜'9�]�_g
��K��z�b̺�@1�W�����h,z�	��L��U�S���i��O���?u��X!��6��%o�K�F��C{gI�S��$���
Ĕ��f�c��z�G�u��b�8�P�8&gME�6V��8��Sn����(,;t�̚��`������l�����|9xwɘ��sZ�N��Oe�7X�Av@����f; �D��wNÙ�c���W��Y��R�Y֧< G	����1o�[��W��^�U��2�c�W5�N��H����-�4�
ٽ��}e�Og,����y[N�\n'n1��]����9u�pof0Qe�A��a���ݪ�.�Nj��͒�"���/�ۮY�҂�F�IXc��.��+9"١d��=�rV���|��OT��k^pf��RO��'�D���zQZT�������*�\��,�[f��;X����v��������@z���F�;As���sr�t��pdU
y�N]�W��T�n�8*$k��E!qk��=�Z�)�pu_��I�P@�B4�x^�<0r=8�]&A�^�h�H<2MWoE��.��p�+A�:��z�[��wT7����NǛ��� iJ5����іϫ��L����LE?{/���@ 5p���J�N}k��9����3Z��ǔ��>�7��T\9v�B+7���'�A½Z�K)�ƺ�Ձ�����K��}��	���$F�}ٰ��9�r��&+�J%s>?��'G�ǖߜv����Bn� 03w���A4�FyIxn�����⌌!�i���?b*�
6�#~��.{M��s���Ox�n�sRcGѬ�'Kc�8���u� ��i8��?6b���F��{ݴ�Y�?�L�D�G���󟽧����<���'1�@oҧ��;ȗE)
wZn���H���<쪎~�-}�Z�6,'����y3NS�W�lb�+ϓ7c��b	n�٫��hx��8�?��kW�[3,e��k�N�F�hH���u{P�s>Z%c��\m�Ð a��5�m
� �T�4+���x��w?l`����q������	������x�.>��H����L���]�k�M<��z�PB<k�"d]������v�g��r���wWq�gi�V"U�{#�l�`�y	���h�r�iըu�mD�
��|��p�K�o���a]HYV5���$������7j��~ɸg�D2����۫pÃ  E`�r�x��E�ؤb�a])G��\�[�����os��Kxy��}��d��/	G��Psf��P�l�6��gkN�`�p�f�/��3�U�t5�^�C�3&?W�9�᧪r���H�$��鮀��6��O��c�DT�o�6���7 �Y�7�x�e8E7�,�z�]���C>���G[��R�#ټ=t��cǸS8�I��О�mO�d���'g.uN���ɏff���c�y@�[!>@þ��rm����o����Wz��&G�Գ���w���4�pUt�$d��x��a?�}���n�2N��Zr޹�	�JD�N��<눣��Jz�C#�2ʝ%E�'o��!a+�����	�4�Ӡ*0ݮ!"�#��˫�,���zv"���nD�?ۥ��I/v�%uo��`�3&��:V��z�b֦?��M#Ai�>QC�Τ�i��ܛ��!�"�Og!��5===p�����A�fAzyaH^����4 ���߻զ����Ls���v��W�_X�,�
�!�~�`g ��xŝǖ���������uaes/-����E����oڏ���>�������혭�[�GĲ^�EN� �do���XZ���`�g,E
��g_�Ɖ�A(|A�FC�`�p��zS2B�,c��;B,��7ćŏy$�H��ٍ&a�`N��፨D�M�F��Kh�U��5O;�t����)�I)X.��k�?�E�fH�{&���~~S��ޕ�S��jE#���:X� �
��
��ӈ"��0������Z*Z�������Ϧ�e�� S��{���lGח��}v� ��]Q΀C�S�7[/Ý=Hx;�Ν�O3���0�_�D�9�e�����x?^,پN`ȅ5ʹL��~x�,H0�{rǝ:�|��-�.��L)��-�����R0���%^����dH�p/&B�ER�q�>8,+0�V,{YX���$����2у����<y�_���� ���@���f#k/i�8o���[^��R^n��T��x��U� �G,s��~���Ƃ��\H�nVѳ�9sƝ䑝��P��oޚ�@��ŷ��m��po��bF-��0�!�\�yQ�ݕSAP�N/:�%q��D�ԟ��1�=/-ؑ�m��8h�����T���68�o�3��3�5�Y��ٔ8�xo�p΃�3��{�ej�1"+���&V
�;8��*«!I%���;��Q7\��)z��4��$}Դ$P���%���~>�6�8-��GT� {5R54�D#f:L�R���3���|%��%��ܹXN��݃ɺ�Qβ+3��(�Юp9@:!g���)��?s��Lq��u���_�Yns����YbPSu�V3����$�ܱ��>����n>6_��<=�0���5���nr���%˖VXk�𮽘��Y����0d����|�B1P�ڤ�@��\C�o7��6D宣
���`,�l=�!����kc÷v겤�+bAis �t;�0j�����2�*)/U�gطJT`
�� �}�7��e!ӌ���T���%��IC>��f1t���o)��q��s�:>��|1������%>fVe�^|���6�T�^z�q�JX;s�ڜm3h,}����
����Zآ u�0�J�U�t��h�v���F��N_�ژ�V�1n��wǖ��6��O��6��5Պ��r���ݓ2�3��d/�hx��b��p�����;o��OTZC���E�P)��CWp���}Yw��S,"yHw����>z�ڗ�g�)����M9�
'���0�����j�]X�-�3�Y6�*Ω��x�@���!K�U��K2*>p��~?VX��l�z�B����cƇ��@Y�z���V9�>�$�E�y�gbXۥ�J)=9AП��iH�Ɗ8��9��u�	c�4�i�
&4����m�(��.%Ŭ�_�3�|IhDC�c�h�������_I�f���
�e9���fR��s?�;	�����]V��MTk�����Z i`Ī��� ]���Z �,�b�3§P]�ɲ9�=珌s��#�o��^�|&�5�*J����I�}K3���+Թ��nB��s�����0�-��u��DT�$��=�Sg��Ӹ�_�_p��
WE��tU@4�pH�;�59�<������<q�sG��Qי�쯯�<���T���F�c�P��U�y;�H�pL���6�n�=��S�ξe�3���o��[e�:$�\&����s�n�^!K�I&/���z<��t��dU��J%�?�йL򨒂��F��B��e��'�z�FQ�f~�ua�z;�5�U�0��`�t�$�����Bݺ��{-Q ;��\ 	��)`ȡW4���Ո��h����A� �Ы���܅PR���l����!�8�E���G�/�jEzC�b��?������9�y����4/���?�Nάs�M��QA�,�����֛g��=�p�ʔ�s�=����p�j�xmI�G�!�*�;`v��!A^�����]� �L���^�w�^m�`*�I"� �ݹpG�i.��Pn�hw�2�b��M'M"-���X��nx�
�-c�`�F�.,P	���� a��m"'
D��Sڪ�Հ�i&����QB�F���:=�Y��/�qű���~j �7�g�����N�`w�7,1��R��[K�x\[^_<�@��JTl�Q�2w�/F�چܿ.�����f�:���q+ls��E��;Y�l�;S��fb"��*��~�h@z�?͞m���a�6k%7��}�N1�c@���	t	֔1h+ʱ�H;��� �"ˉ,���o���$E�]S@�&�1�������{xc���.kz��1	b_t�Gu�	�>ob��q!�4V�Z����w��0^d/�TFAeͷN�F��c�iW���݋�$r�Oxh�l7@��	>�,
O���w��ȥ��kXy3�s9�v�	�~������R�8�J��C�M�-{ȝ����E�������yO��K�Re]��wm�+@4��A��:{�;ϟ���>��-d���v*ja]��TvY&n�_���W���wi{�f,�Zj�x��\E�z� 
�x���<0�ms�4�ڨu�]L�é�v=97�N�pXN��#� gv�'�?.sw�Zߕ��T�ADau��ޞTVb����]�h'��5]Oڨ�p�Q��o��7㌒X��c��ϙ��WwK��hr�(_8%��B�bl�S�z�s�]�`��^�.���۲���t���{=#��1m���Ŷ��r/��zC�-����k�>�J��&�-z2K��z���^n�i㪀�;�o0}e�%�W���R��yB��1��Ub"��[��Fx-\����/��`�ܻ�#7oq�W��[�:�q����YP^���rU�6de�0����T�-��9>�$� ��G?ز�7t�IL(8(k�"ظ�����{�Dc��R�\�j�*��>^"�
8m�l�M�Wm�%� 5d�6m����Հ��S���On�>�=e��:�_�w�!��Ms�[����=c4X�a'�-?���FJL�&vC1��9��8BW?�)��J}�_o�NG]C����J�DN�NdY�#XlxV16EB    fa00    18a0����H�%���V�dt ��1}�ҳR2㟹��$������[��M��h6��$��Ɔ��]^�d�WY�_�I��+E�n?�$)z��>@�S��ٲ��m����u=ūm,j-����i�t�<Z xT̠��h���^v~�G���;�O����s��<;�b�@T��?`��=G&)xa�|���:A�{Q>�*�F�]��0Fz�<F	�����=�r���C��~�EI)uC���r�4��7%b�H�+H�`��(�uDdA��.�<�Хnގ�|�B5�Ec��1�2�Y
�HLc�߈���Iq"tqEm!F�6���3:0j�5��A�v5Q���P��[�}��b��zB�bx�ꓺ�cT�|y�����a�:�Wk�������׸1����x+� �J=u��u�h����G��� �$�Nm�������A.˸�h{{�]%�ָ"1V�4:�\9BS�iU�-����5246A���'V�p�.��'?w�Q �^�i�*wEU@b�:�՛u��L*��տ��l8������Ũ���vj���9��G�L�}���^��̨�`k0����k���6R5��$�@�nr�a�o�y����7i@3v���Y��Jwm�*3�4���ㄝ�C��E�ފ_8��y{�]��J����@.�Da�1K1~��PB�μ��s�5�&i$ x����D+�\:���4%����
_Z�0��O��γ��Y���Fh����6���*��=����������w�H�O��s� �}~�|���[�^�q��.���A��(D��AM�+��u'�U��3ׄ�p��d�.(*�~2�fD�a�_��1�eމ�#[��<���at�c�V��i�'1%ӑ���!q�����+��"�	�+9[��֥?���f��g�%�ߟ�>��`�a8=�^�Ł��i��&�y�kn�ʼz_gƞꑃ�V�I���t��-�U����͚F����kL��a�W_Ɔi@�ڃ�vpC�KF2z�bT~Q���(���g¬��֑�������	Zm_����ߝ6F��ůȿ5��O�y�4�ݍ� o*[.��*��ҫ�q�߰�W��G2� S��%��.;~~�*����|<���<���2�7}ǊJJ=돫-�=���ݾ��|��H��Q�0�T-���갅��rF	,�T:���.1���A3l�=� ���+n*$��v���>�
��<�N'���a�:N<{L�`& }FD0�ŝٔ�t�H�P6��0zx>��5���/�_�˺��IRS<۝y�x"�ԉ����E(����6coY���m���L׫�h��}�K����ؒ%N�~��y$�+�..�n��t;L~��k�웠����C��E��r��K�'	~��;�F׮r�/�?�ƆP��V9�7�N^k
R?e$�Ź�w�C����1pH�I����c��5�þ�\a��H��@��1���� ܵ%�L�:�|)�n�!��l���'���?�g�Z3�Ox�g��f��)U�0�-R�̖�O��;�r���w�-<��"�i;������*�T���i�MG�P�Hڌ�1�~�=��x=�{�Z�m�ӊ�C����o�R�T�.=M�V�C�-��ϗ'����%���8��&��mM�F�������]ε�~$�b�>����I��� "޵WVR��b�;��Q��q����Ig�bu�G�a-� X��L��)\k�� 	�~�܄�C������MęI�YY���V��D7Ǚ[����Q��:��m���R1���Zz��疻��W{ZT���2�;���3\֊�Y�v��YL�Н�C�M���<a���o�;O�=�sJ���l�^�~�إD��bM���p��ngQܒ�q��FI<p6W��P��S^,"�N��8ȼ�2(r2���`S��O�0���FK�_| ��J����Y��V�U��5�!�8_DH6�˫S"9��4u^���:����l�l��}�ǚ�3#p�{%�T��Xg׺��l;���Pj��̺%`Û/l���b�A�w��:å�r�S��2k�Av��]C#�RɒQ��ĽNY�u/e؛�<�����x�:���(��).�/����d����L��;@��`�մD!����Aa�ys&��)��{�o�q0����0��d@ ���!~D��L�`�;�1.��'�Cq:�fVQ֙}_�9��B�LP��Qt�w�p���7��o�bn1OnƮ�� r������?B���Aq�������˞�Z��^��2x.��u��a�:/�o��p6���@��,�,SG��82���_SZ���p��T�qL������E�8_S	#]e��=�#-���,r1�8[��7`�hC�٤�l>�]�}�-<�BS?��d�ȯ��hi�2�Wd_ 7�a�,��ꎺr�w��(ؼ��*���fW�dg���@����k��Ү��Ӱmw�/8c��"��i�@�yV�OΊ�V�+"|9щ�(�D�I���;�֖3���������7��a�e��E���Y�u�{��L㔣d>��p�7�a�[���"��K�jǃ	^���?�Q�	.�MR���U��Wc����b��F]��{EP.Ƙn��u��$68��g2��6�$����9���@���r��O�����w��e*Q�2u�| ��r�t�C��5?ē%uo8�+�LJ��.7y+AfC�����r��\�0�%>�]��{rv�{7��G�d/n��[�5���f`S=�������h����|��r���?��&p�s�oڎ��Ҧ
t{��j#�Qa���f�a�r|E�l���A�aZhٴ�����	�(��J�y�|��H�����F�5�|�t�（>#t*R8�Л�˩(��(��Y�L���� ��s1���4����,R�⋦oKđ��J�2�>��'=N����e�ۯk/�ߪ�?a��Cx((O ,�[��N�S�`g�C�u9��N�T�o����k.�n������Ÿ��l�f�l�o��S�a����_q5�����꟪���U�y	_r6;:@��u&�3���{�˦���.׭�n�1�� �R�v��?�����]������?�Ų��!+?q�PL�"dn�9�|��7YK�+u����B�[7��S�g��AG�SU���'U����D�t"r�E�5���;ޯ�`�Ip��0�i�7��S���4T"�]&u2���@,Hk|�K�~^����џ�o�I��s']�W��o�!W[xWn��Ȑ�m���$E�_5�RA{���)7Ȁ��Ѓ5=��c��U���DYu�p�6���@�P��0��
 '�����#݀"�n%a�S)���k�x+*�E���a@#����b(��\�U3��k��ﰼ=@%�{`Mb*��|xu���b���ƺI���z��!�0��q0��*!��$�n�.��k��[��� J�6�L�F쐴 �b�}�H��;l.Q��<	��96�?s~ݮr(J�a������rw�*MA~ �Ēj8U) �~T�����1�%"�A�PD�,袁M`Tdi3�r�D=$��p:Þ�L�������u��f�О,��5��0+�����%��V���&�]�Ya\�d�W0��@,���ꍎ�m[��{�"l'�|���� �zWބ���y�X�ugj�����T*����9�1�P�M8�y�Z�{ŖXj�*�,n�e������ӭ�2�i0�:��a�DA��h��^w�9��������ʾ�}��H��ַ�Z7�9�9�\���Am��}���S���:
�]��f���O��/�'�J`����UM'�1��u`��W@����0��ï�š����q�����kn��0��[Dʍ��ӛ�c���0�0�U{�uQ���H]�؊�W�y�:��;J(R��)�_a��a���q�H5EF�kpe� ��dPRS"je��pW��Y�L��0k%�eF��&�*LǄ�ymή��n1��S^�^w���S�c�3���}ۦ98$[�/vȥT�mI�p�x�� vx.*ř�"�n����k�m�_.í�N�v�[�yu�d<�����E��N3i�g�Z��i�Ȁc��ej��S�������dd�3±+���ڸi@����r� I �}��͞�u�`��}�v��x�J��P��f0����ŭ�ee�TT�S祂?[-$�I�%n�,��~��^�S�
5���}#w� �d=��N)3P~�����W���(��x����h�%�R��^cE����b-�xD��GՍ���B>*ޙPg#+Z�
,`��������,��Ev�"v-B��5�I��N����J��*#�_a�k&wP���a)� �l8���@++��S:Q�&C~9�Q��V�:��E^�kC��[I=}'��
�%�Ӹ��=V�	1O,���	9d�	��e����z�LY��uD
��#��m�lg��[�t�լѱե�e <-ظ�+�Y�9�ט9�+VV�g�7����I��z��/��/iY�W޼������$:��T�3$,��������X�C�Ys��/bn����/�3ڽJhg�%al�������5M甚r�r%�.r�_Z���ݣd[�]�Ӯ�ĝ�cZ����G�-��ұ�Q��Ji���˴�¦Q���I�N�������\"|M\��)�"�4��S���DO��%<@ɘ�^CL9�(:N�9��8�Q�?F�'�N�a�F��e���(��6��h��Z��X��Y�b�)��~ϯ��˺f��:"pa�>��G��b�~�����<�������#Q��G���K�{��P�yF+<��Ҫ�mt@� Ĥ�&����V>4��^K��f͑�q��R�����|GJ��H�A��=�Hf(�� �<ܦ����sFv2�~�q�������D�i�C����p�ȑ������ϼcwK2�ɍ���
�{�-2&�qckw}(g~EL�>�6��[g���u���-+� -y�����'��"�'�/p$�^Ԥ�0j[�y��Y�VtT`��b0uP���D/ۿ��4���8"S�<�|fKӋ�l9ȋ3��S(x�U��6���j�+2c���m�7�ԏ�r ���˚��I�I)�Kl��F�Ӽ頞)���rɯ�����c߅��v��3��R}Fp>���O��)Tz�� }�!G2�HZ�<�"K)�'�� 	f>�<�b�!���V=C���»�����kL�5T�Z]�)�ѕj���4�J��t�u�}PD,:	m;!��-�x�!(�����(���2���Aի���=x��Q^)_��)��:�*���;�أ}�K�=P��Z���O�wKx��wz暿o�,^��>Pk����u��+�1�c�ǟ�&ǹ��Onj�x��І�յ�V��?򃍁�|��u���c�B"���	Y�� G�����K������uy��ǊEM���A��v�D5�g�g?aכ�&��!g�K�<�⦿\F�0���	��e�cN}���ø�����7v�9�F������Ŋ��^Js� ��ɝ��OW�T~`
�£�kT*�i�FA��Ko���3�<D�~܊o:,	��VMj*7�9P P9��������[B�ڴ��)֍�#��݊�D%7����^�`&�d^�:P!(�tP��+	�|�x��Wi�?Q�f[�LOL�������I���A��0����Pz(G�|��灉�I������L.��uY�r9x���/���D�We���P������M�������T)�� %*� �@�x��-H�.	
�"CZ��:Q������'<�_E�(�[��>Qހ�m�m�*���F]�/�`�����'!��Bg�R6����4S�p��?2i&�q/��dup���~�Q�R�g^
mSy�z��F���ix-DfX��^[	;C���\T�� �s�#�qX�Jf:���|p͐�+R�yK�jz!�z�΃� �B��*�����&7
d,�4Kg�����ٟ�h�MU��l��^�.�v �}����c�d��/�ڟ�zT�����(�<�l�XlxV16EB    fa00    1a20F�/����S�V�bV`�h>�]H��@.�4��?p��0�fP^�pD~�o��cqy�~`��m�j�&R�I�V��dQ�pX����j�{O򃁈U��/x8+���.u��3X�k���/�P��d���^
��wsV�+;x�2���@�]��v,�^|�Md&��c�ݯf�X�_�h�8A�q��(�Q؆Ex��Q>���|bRV�d#�R�BWC�8=�֠����9��Q}��4�85<�j����ɍ&���۶�&Ó+� ���@,�7=�ny0�0�,�Hr��6U�ŏ���̜Y�.�z��E��gn`���û���'�l��R4�����4>�Jߔ��o��6=/�f%�K�!$�_"�V���n[�4�U~�`c�#��P�M��3S�P��a���t��Y�Պ/l��s�K�O�qi�m<�6��<t��ș��,'y�PnYR}W� �W��4R4_)����؉�U�ݱ�}@KF%RDB���R~r*�#o���\�@ִN��_��#;x�
�*�H�%Ѫ��A��;@2}c���_�]�gL@��(�ե�3:9�9[桽���y>1����0/��3�
������Wd�L�I1(�������vV;�3S��;�צP.��T�^�s+i~�$���G-�k*26ˤ�.N�����<�N�����sC���,>w��O0�D����l������w�a�+�?���-In�0;��6��4l�n� ���CSX�|w�]�dۡ�_�M���4��1x��TT���޵xMO�6�G
�4&�g4��p�T����@�a��o-�S%��"8�1�5.�'��<5��W.Y�m�bX�ʻ��DMQ�觭��>i���V&	��ÒWД0kF�-��N��D������n[�j��F�p�� Lb��]),d3E�U����O8�(П̿~Y��p�_~].�`{��~��lb�d�ڏ=�Q�6՗bt��2E�K�cD���2�Z���ZC�u������f�y�d�fL��G�����H���ѭ�	|�NL?g�����H�Ix ��R���U����?��D��I�����=�١{h�љgEY犑��j�¾������/	:+�!���1u����`Ly" �����A\f�t���,|���xW��b�;�
HI��a�)������m�`\?m�D�#�+ra����h�yB�A�:�I�9�d?��XQ�anhuk��������j8�Í�w�x��S�d��q�SLS���]��sS�������S湿6�Y��7����Vb(��1<'����}���IBB��}�Tua�n!+���<i��g;xT�8ĺ�a}z����/~)I�"j��Xk�j~O̗!�X d��ai�F
eDI�x�X����Z��4��6E1���y�nk��*��	f��@�!���V���?.�!��g��sW��cN��B��kO�W��U�H�D�%��-��O%&>2�i,	q��%R�lG����d�GTeJ߼Z�I�a'��u������_Jf������6rxxĐOA:�_�_@6&��%�wՐxO�lKf��Ϩk^�On��n�A�˽g��<���6j4�vY�
��ZT�/`~��y��.��ȣ峤����RE=���e�ے����r	*5��7��Q��<q=s�&�k����M��>�I�f�:��EŻvwa,��Ux��Ma�X��*����F
8����ԡ�"T�@���g������?c
?�WvJ�&�n2�dy��_���B��uLf�By��H�)e�\�K��h�EX_���1�d��B�j[[%����!mϹU	�R���I*�	7���6
}-7H�O|a����u�켵9���8}�#?��{U���(v�"�����F2" �o^c�'k^f'U<��t�Nl
��>�����������c8�T�C�����]�D��N����'��v�ê����طɱ��1�4� ϴ��
�>4-F�$��O!�>L���c.�����+����~��&�8�N��w"�$���L�Šܒ�2*��I�r9f�B�晟�1'A�4\����C��xP���&<"S���[��J �����"Q$�h�4�kV�-�?\���v������ݯ��/��v�D�M7/�w6��]��?S�ihh�<�2#4h��N�].�U�f[�xN�Ҫ-�n(�<��Mvʥ_�<rbA�?�(r�nV���ޱ�U�>���{��kJW��ӥr�z4t�}	UqE,G{�%tJ�����y��+ՀƬ�5#�j��4K�v#G��n�;������]��r�%�=��6S���0X$]��Bh�o4��Ȏa���x��a��Q�Z7�a����*v#����y��ԟ������L�⮂PKV.�4<���ܤ��j���&~o���T�u���I�͏G�p$Ȅ\���}�n.����n~��6���3��u�lB
���$}<<+��M��Я��0 }E�(�/�ԬG���L������������h��t�?�p�$��t�hMqn�`>Z+W�v�k��]]���N���E��!�MA����/�$�V�8D�l��L��Y�g��+B�����h�b@H,R��V�!eA[n=�-4z"QX8}뤐
Yz�bE�c�_/h�#�U���C'����䰝�֗(1������	���C�H��X�Ƒ��]�7���Xl�	�{��m����-����Tja��9�+,�@i����z(��,A;	����{���5��R�`�V���������#�K��n�hA]�嚴  ���ݕQմ(��/Rd���슕.(�v��g�3m�h~�~=8��n�Y��с�u�w?%>�AbnG`��8��yQ!!����f �z	J�:��u�鯞A�(�[~����KK"�@Fl��:&�$�~�������]5�?������Rm�1R&��{��n:�<h��Be��X���n$��yQ��2-�OJW�[d��~�����VB���M���MW�(��"����L���^��S
^a���_^S�A%���y)
$�F#�l1|~�)�����g�����*rj�	�ˡ��-�_>1��0�l�~�enXT�u���l�_��O��]�B�v2-}�m��몵{��x������|3�����Z/���D��p�Yq�ףy]o*Z����4-ݚ��F�e�٠�?2��^���Ҍ���q���~�[�
����	ۓJϫ����cw��j_���Э��;�asp4�g��	��^��=qd6l���5�-�E:dz/x��(v��B��򑻧b�C�.��Q'�!�:�y���`ӟ���p'�;�5Ӯs�`�Z��>��6�aNV#�o�����BFɪ�J���U�p��^~��lx�:�Xp��%S-�T�����K�C/RE;C�%ړ�ʮ0"To�(on̚���_����jR�	��7<�s�F��6l��El�����^�,3*2<�N�|�ҷ*�:"��NT�*�xƌ���מ���瞮��ή#B���1�(�#!��=*2�N�=��>
W>S5��᪰�lDY��S��������n�D)+atFPa��;fy��zR�>N�W�]����lTU,�\���0��y_F#�Ě'?P�UF�O�lL"�r
rnq�-]e�䵩�����4K����{�Z������ٱn�w߫�"�r�f��o	x�YI��A?��9�/d�����/	�n�R���� ���7�P#zdu)R�{[Ǵ�`]\C�&�Y?�Μu�Jf�"r��!�d�=�X��e�Ǉ<����V>��-t:��P�碯��I�d1�XޡR1)�����!@��I���sApybԒ�7�Z�I~��`Qi�7�lq���MdZ(�y�w	pO�
��Y! I��_�'���_������d�ѣ铋J��B���<?�4o�j�����F�
?��v��B��o�m�����0yi{�&��b�L-�Ɠ�
gS���?O�o�1��u�zp�@�H���)n��0t��-�gA�|"�N��2�ߐ���@l�a�� *�5�K�����M�ACf^��f�,=��Y�i��F_�������T�m�2)a��F�.��.�Y�9Dj��>�j�jT���c��4���֩��v�	�|#�J`�>��W)�q��C7�1{� �D��1M����ᴸ��਱�54�EߣY�5c\���wI��c��
zV2�j2v���l� ��3��nĔ�.���2�O�O��(����8X3�n+a��"X�>q�9��ob=EL�$�R��*���'�7<�I=,�U��f��T��5<-jS�n"�W�6�ځ�Z�ݛ�/�ڗ%0�w>��l�<lƆΏ`�*��Bj&���@��ʽ�ʂ �u!=���5�f�[���D�@F���h�y�[���3[��x���=<�dZ�J�h�����a~c�Y��S<�z�k�D���kJ�5�a��Ǧ�)لwJ�\�6z�Jn�ɒ$*�@���&ioZ�oB�A�����̒`�����	�A�ĝd r��K�S��6������볦m��`JѠ�ܫ��p����K�r�'�W�Uy��]꧈&��!��\��W��plz���*7�v�W����޵O�&�]�r�����7���1Xb �Q�
��0�|:u4�>7a$]V<;�MZWd!0�Ȳ|B"��+ n�%��[�wnKW?E������B�EhKY�J�;MƄ�'X�)���b�7qʭ�"^��|�:�YN�/�P=�+�5��o���g�%�`%c��`]X�<�(cS��R_т�.����t��
�\����a_Z`(o	Ȥ�.���}�j��9͋�m����-��W�X���1��A�a�H3r��9���5{�AB���M��Z��� CU���go�aE
z������!�dm�w�J6��@l���>ZZ�rQa��;����h��8حvlͬrf��R٠9�A��?:p���,Z�Dmګ�{�1-#L*��p��U�� ;�nKe
 �GVgt�e�����*)�� 'W%�F��R��3SL�9�r�x\��t�A&& ��fZZA��+kJ�i�=apu��
H�6���n�-\�DF���~�ĺ��2C�C�Or�����w��tB�M�Y����6PSJQ���IJW�-H��O��yȨ��F5����hs���l!=��7�I��*|�\@��>~��Hlh[\$5f�Kf��N�QQ��.�f��2��Sb���c5Tt��vzG�E�\�$���{��� ?�����ݩ����F7(9X8ײk�(F�'N%I�9�`�U%���d��ϋo�m.g�?�����fbL���]���;��kY�B5���S��o�ǎ�o�Y�����$�Yw����TB ��>�����h�/g�{;��� @]c�8?���7}��!�E���FSc₺��3�1����'X���}IB��4[�=A�C�Ápo#������ ����V��G�C�Q�g����z��s�T���W�.$��0�}f`�|a���Y���{ξH�͉O7��PE�$B�	�/�p�0]�;	��[f�?���	
Hh�.� �G�����ڀQB�a	��6|)�B����ݸui�ڳ�}��3P��:n�U�t-�#�LZ,��X���V&N��7kčw�V}~�8��Z���xY"\�qJ6���=��^�ԉQԱ=c3�f`�-us��:o��[>���M�.֕����/�_�!����6b���]ш�O������@hU,Iѣ�9`��V$�<����}��Q��2���}��Q����vD%Ը͐$�S�8��b~���`�N14�V/�|' �j?�g��p�/����Ⱥ��"/J��mt��_ѻ�9�o_��Ԃ3�zQ�p��%(!sn+�E��}npB��;e�
�n\�tUSS.������hM09���]A�Rg�
��{,4-�"1�$�Tّ��iw���i&B�>��f��XL`����&���)e ��R���;�i�I�>w;ekP���Q���ж�X�Ylv�Sv��?Qޛt�=D-�ބ��&���9�s�X���qq7?�$�%r�1�4-r7KѧA�����^����$V�a{đ�-�?!Pɵ�}Û�P78��6�z-u.I��R�>Y%���S�_��Vd=M`%v�Q�zd�9�)�tz&=�?���;�p�Ҩ��w5I7�8�h?�Rߋ�z���E�����r:����7����`w�cbɽ�K�y���q�P� ���)�M�v��^�4�lg0��yHc�����<�#ۤ��_y�p��q/-�5�mY,*$�x�uQ��d�P��d#�?�'�g�|��)�|��ૠ�c~z?��n�:�x���l��z�����Q���\�rfj��%i����NEK�|����{|d�E����k%���2�;�륶s;|kQEg{�-!�6�j`asY*g_rl���%cvu����Tl���/�O�	�h�D0��	E#�6XlxV16EB    fa00    1fe0�2w��;������ifv?M�u	������P�e�,�MvoB���) �*|k���������*��/t�J�a�t��O��}�O2�ß��6H_�vD��mq�̈��p��z{�
��j4��CM:Z�B��jS��y��c�o�T��J��[eC�D�]���d
�P>~����tbiǇcy�4�ת����{��ª�<��f��-��\c�q�j�c��JJ1��XP�]2���5�"vzy~}e�_�!�h�q����}�Q�і�����	.i���äV���|'���_���}&I�~�~y�3`I?�~|X$b�ca�Խ�.wo����sb�G����YZ�֝���A1�AT߀� ����X�/q���v |�Cc+�)%x�� ��6���:��\��������[q��6�q�b�R��&=��ɞ��(�b𐋽s{d������Y��b�A{ڌQk1\��zc��BB^�>������ݟ�?�����-B��oۆ�'�5��.��� �|49�y>�-|��m��@#����5mu�$�C�5ς�}��<�^=�~�':�{>��V����ࣨ��X��S�˒��1u�����,�ͧh�*�m*aI�n^)��g���BqMcOx������P�G�Ԙ���	dD}t
T��<�J-=C�%��7��/�K,Ն0"h�}�p4]�I� r ?��K��%�Bq�,j�M��gt�ǐ���]���N��:�6�܍�t��(d10du�kTt�ٔ\�a��X��.���Y�'���-�{l�N�M���c����軟T��"��
��_r���Y�z���a3 ���J�Ur+X�\	��(5�}�K���݈�0�[G�ft�z�9��C���r��z���n��)����i=D3�E�L#ݔ)�����-t��<�D���,�K�T|��n L���׋�1��P��tnQB5��˃L��W���R'�̉�����s=#��dg���sb�^x���M	wP�20��%��0�_˞&��������"9ș����0���x�Ԅ���sb�WZF?�A�Ԕ���EL܌I�����p��V�4O����{k�{��]�H��D8�~�+�Ҧj��5�nG���>TsX�M��E2^vs9���I$D��G�m�	L�R���@{evY̵�������&%�=�����e$��y�u�+k���3����"?Ъ��;xA��jI���;i�8��6�o���C������VVh3`a�Q��b�W�N�[9�[s6�pN�31��,k"�z�󷒞�]��5�UROyϽ1��}D��L?�� ���9�sލ��!e��v)�,��hWE�I?�L���Gv�D�����Z�Ϊ(�+|%���7�!��B�j�[�5-�㩦�w
�,6CD�C��m�aI�~���ѱ�?n��\Z�U�N�x�BD�BOA:4�Z]����r
 ,�٧��'j]f�e�ȅ��Oc�	Z��^�ӊ���X��0u�f��gI��KxmԘ�)V7Jc���>:
����S9ש�c���;ʆU�g�Β�wd�i+�T6TV]!e:���?��/9��wd}�Zz��8�I��Anq�w�]���#��\y��ewtO]��5�o"��S]@}�Gǉ��:��"ª��u�C���p�ShCl:ŝMs�Y�^R1�iӯ�[O��s�	���X6���h��w�c�� �v�Mmg4n"�_0��ѻDC�A� ��7;G�T�+������L_�J8\��x�#^�V�k36ݖ=Z!�f�x_X�A��z�(B�E_�+���{��(�Ŀ(��f��!���g��U;î��Vw�ݗ����SwW�i7hu��ܥ����I�rH��?R5J})�Fα��u!�H�x����Zw '��&��o,���~������BŲ���_F�y��J�Q���B�P��^����V�b}���S��P/v)�#�I����v���.�}�GвTT������h�0}��"�pH	�c�I��!l	/!b�łS��J�x ����2�ڶ��z��cu{��ai��.O 찰tAcT:�R�5�3,j0�����q�G�--}�8�b���7P	ײ&�}8q	$�載ȴkv�(���';�X*bV	�5G��>95��L�Y��(�� ,���;'u]*\� �B�����w�APS�}�/�7�4q��ޕ�¸������x����ű�IF�n��T�=�Mԣ$e�L�+�&����ߺ�S��cڻ��cf��l<�g�D"��l;���K"���s�k�Y�y�F�E����l�,c�Ԯ�Ӝ�k3��vKn��D1�S��{������n��|��G����6�L^�t�|{P�w]:���6�t=��	s�+s�_��ja<�K�����u	�x�q�dذt��
"����4��$�v/�O�V,il@ٌ������ai̊�7��@�a���&�8G���f\z~ˢ1�5�z��A�F\��J�ݮ�O�w�����8D���.V��c^��T��%���F'ɸ�����=��TF�	[,O܄�!D7#���kvc�4���E�(o @���H%:b�ɓ0�q�O|O
"�Y�Þ_��cv&�?�y���Q�&4a\ApHh\N�!��|�౵ĎiY�n�/:���?󑯃�Cˤ�O��xW��V�ZӏD;��)|��Mv�x�J#���L��W���M�;�J��N`I/�5�B����`f������K[��P;/a0H+���Tا��e���=���-"��t�{~��Ͳ�1-��do�`w:nk�럴+¯��µ�=��W-�^�1��*b7 w���Ϙ�;����7D����L�$�!6o����5�*I9��O��~*Z0.*98~��}�|���Wy�������Q�4z�z�nf\G`���\��O�����u���Ǣ���T��{�(������h�.��� U�L�&H��H�\H�=;` X^2��$i�aH`�+�n�J�v2�R���5H�i�!���A�N|���+:�� a���~��llOP���ڄ�M�\�T?�����A0�ĳ�7^��,�s�ޤ�e̊���z�����o�!�;/<�F�MYA�!�)��5�֊���Va���ҹ�7��)��I�<^�b
a�1���͌+�%x�_W!�Y���j]X!E�m4A�4��I�<Y�׹�o��BF4ڄ��V ��"���0T�V�oY�P�:Pcޢ�9�A�-�I#��4�Գ5w_r�}����9��jv �?W�?�1�Yna�e.L��=(}�H�gNZ(I-P��Nb �}>~V�L��ŋ�9��5��/�z�F��Ha�d�|��ß�$T�����b��,���|��7�D_����.�"�4ժ�-�CѺM�d=U���8dĠ<W4�O���o<9,}mY7�b5#<AZ��Y�X����t�6�΀dyw�+���J�߯���w���s�.�i.���_�FU���&�G޴�h����pM���|*l�������ht��0;�J&h�V݈l'v,̢�H	�=��y_�oL�<	�cD�M`�Y�<�U�è`V�3g��o��طé�m�Z$��ad���2g�ё���:S�z���]�d 6�j*��&~C���S�<��4!�@�:�I<SG[��GVWhq�0��.�զc̝|����by��Q���P��V�ҩ�{{g�y0nǾ��h�#m�ܽ*�����k�ρ��NwPѥ5�_{{x5#�u�N�~���}�x��X$��-;%?k����[�J�)���5ɞ�v'�m�u�M�� �+5Ǒ ^P]�C[�47��ʥ���[�<�s����/1����S��,F"%P�l;��\ ���̿��w-�v=��� u�ـ��ؙ��������3�h\C�u�̓�
^]���[�!h_���H8��J�$I����-��U�����т�J�c�V���R�E���j�P-m}2�ٞ�TL��|Z���8?�l2~�A�AU2��tXV%3�è�?�����W�e��}�X�Ҫ4!'&�)��1��W�u>:-��@�k5���ě?�G��@�%��`,��.
}�jvB���&��������~���'��1�Y���6

�Iz"A8��	�r�� �PL!�����X:�fM�K�Bg~���NF�0���%��2����^z����uʦ�{�n�O΢�3�κ�L�eZכ�Ƴ��-�<D7J&3�s��/���M^�Q�0-�q�Jw0�?�vX��Yi�7�1E�+�f��q~B)��:�������!�����ۛUY�� 9u{$� ��H}��jQ�]=�f7.�g��<a5��K����yK�V>�E�D��f#\���Eg�!/ �@�}���p+���$$r��d���=6�΂�^�{M�O�ɤ�C�Ĺ�6E`O9�}m�9�v(̕?�JG �~T첟H��ְ0L��WR��<��&$w���N1�q�W�[7#:�./Q�'6Z�A�J�Ic/�����^��(=ɒ9�Yj�3�P�p_mJ��A0(��Qdyp~��߹�,�>�}P�iZ�<p�w*�x���(�Kړz�-.i1j�C��2z����Y�a#��-"[�y�W�*�e��|,�^�,bl��?8�H�#`�1+i�z���ә�`^�߇@{��*1V���^��ռ�Bm�r��(&��@�[j�۾�X�:6�;�IT� ��SV��l�"+d�lZF�B�A��!>K!g�"����.\	F�?�\eq�$ӡgq�nQ���d2�2���h�HͶ��ہ��7M�z��$�Pz7��!�B��U��	#�֤�'"��Z��Kز�$�#ަN��Ďp�L�H��2�%�汻��on8?Ñэ=�	�۽�W�Ȳ�����u3�y���u ����4ӆ=UΜ\D�U��2��إ�Hɀ�
���] vF+0��9+�t�w3���'u8Ȫ�j1�R���W�ڟ�U���@'���鷁d^��3<x���������'v��(�Q��ճ����E�����ic��
����H�^�߹挩O��cV��v�j &�Ѯʡ��[��M���N7�R��p[��Ģ�5���%�28 ��J�d�(�3��
X7���[z�+�"���a�$�X�-�)Se��vȼ�S�db���Q������er�������F0�!6Lz�u��毑0X�.��J=�M��ys�;�@L<��j*�&_���7��`|�	<E�w�Ֆ�-��F�|7�Qy�ڔׇjV7�k<ݣ�*��?Õ�P���U�&V��GP��˝0`�=S����t0�ޙ|������L�
�q����2�������s����*�d�ۀp�X}���E�T�cɂ���W�*%e4bɣ��6���ْ�'?p�Ax#��ϮL:�T�c
��:0o*���ƥ�����j];��P���RPA#��B{Q�����$ �}i��9&�&��%��3�����^L Td�˯t�iv9)�����{|pd�K���K�H��$���^��uY⏒��8:�WUs�j+d&ES�%*��d��p�o��Fdñ x�N*���~�EO�&h�(vɞX�&�L]���-�V!o�&�i�S����?���~�Pl�����FaP,u�$o��_0�����x�:�I�WLC�Z!d��7��ܙ�bW�k�A|�?�g]���2| �d�ݞ�v���>�: ���������ڡW"��A:L�sC1TO�P���A���9=Na�P�5�����]лZX�ʪϥ�{���6Yn�A�|~�Ϫb&�Y�84���x��w=�eC��������T�`G*h;(l������n��fjN#��d�>n��:�~��ة�1��T[��K�?Ӧ��|ZQ�����ss�p��������b��U�2�TY����ѻ�� ��ҽ%8d��o{PՆ���$6�q����Ţ���s��2�Wl��ez%a�s߫��O;�c+ұ��S���ګ�ڲ���}e�ҳ��bw���jT���"�A��$���k[
�͖�	8Y���l�l�O��i��_g���u��q(��2*,){-/y�ʅ^�gkI�Ip�aY/s����YpqU��aø�H��"X��eiVk<�"f��qKw��4�/�vC�f[o?Τ�('�@�*\B�.Ǽ0�g����7
�A��F��$� ��c�S&M�%��9�L�Ps��V��Pn�s̍	����c�`~�[�f��|��3���:\"q-L\��#�^*#Ʊ`�j�bNU%�؝D���N�7O,-Я����j-�AD����<Ao�0���S6�n*d?R����E\��� %5tZ���b����s+����<�[��Q��A�ps����B��0�?f�����N���1�*a}�{�kF�o��CT�}�}\4$1��4�b�D����SE#���n)���hh;�e�Sc1�Ծ��"�i�P՜�1&�ȯt.6�� E�<�.�K�P�Ϥ�PYh�q$���E�Ȍ���'�'i7�bh��EGs^S�ɍ+�*|3�,����"����4m�R���eU�\귟��E�/�L�k��>u ˱�|�4c�� �����˫g��x$V��S�d�"=�1M�!�Y�����%���j�3��i)n���NIY�D%c��W:���蘮ڢ`7dH�V�5|G ΉW9�����a�׽��H2���T���\Ȭ�����EX<޳o�#�>y�~����!mIB�;l���O����@m� uѪ��T&��L7Ȥ�~��*t=qz�f�.W�����f������`c=�
?�p�Xfa�v~nHR��p�G�[��M��g�̒�[�L,����~Q2T��KIF���_��@�ѷ8_�w�3�iD���n+,`U�.!Rp��!�ƫB_���v[�X��-�$��6��=+B�p:�J���d��z����Uɭ&�GŲб��ˈ���XU�͔�r22�X�Wj�������Mm�����G��#�Rn��f�?~�J�<c��m����v�:RV���X�Ż7�,X���"�j"1�i��:82��$��v[t([�%ʊ����|<a!H��D*�{���˗P6!�2���eE1�i(��[���(��n�c�b�ؓ�U���ԅ��|f	b� ���I�Kq.���Q��d��vH~�T��,��c�S�9�kX.>U���ύ"�,gοxn�z�����ÐI��r�I�f��g�@��o�I��m���x7+�A���|O�֡�L��i�x����E@EO�"�r�v"�o��j�z3j�C"6�G��0�w��E��Œ�����|�K����p1���J!�#[����p���J�Vʤz�R��T��8��¸@R%�R8BM��R���	�1��9�m�d0w�C�o�)�4�xE��RY��
�D;��kE"!T��,$(r�<�΂�3�~gPD�����-�̘�2�'7>�b��,6X�K�G�.j/��v��h�z�(�S�4I�����g]Cc��=ڦ�����ȵ-�� s�ޔ�u���4K���-�jBl��z��됨��2����m�?F�=\f/5C����0_�E�~\�;�}���
{z2�����c7�`�mp��3�s�p����b��OĠh���%Ֆ��T�+=V��4j��quxN�����@�+e>R���5��,t�j�3l�9Mm{q�^��9#�p'�t�L�t W��F����t��uNu�Г,���	����~[����G(#q�C�Ͳ|�; ������e�'b�Ssu3�YO���]�IF� 愀��ߑ���{U�łx����B�n��B*�V����TPZW>!J��x�>*�WU�n2�l�3�瓒!%R���ѣ��#��xv�Qbm�dVd���a�i���hcn��2�`���)���W)ͱ<1��!��-5Qq�����QN@��+!�Gٻ(�2Ώ ��;��*����b��k��٤$v�l�H�Ɉ�^P�W4���vT����9�E�'�c�O�{�^�V��#G6��	�Z��XlxV16EB    fa00    1a40�%b������n����gm;^�J
�28��-�5-|`�v�^��VO�J3m��8~��)Z|!`Gx�ݡo)WM�4կ�V58
��j�.=���)+��`�18���1e`vS���TPV��`�jL��r��%.~�t?c�)ӕ�	�!�w]�[�1}�l�<5�y���}R��P0��PO�`��oc�G��'�J��h��2�`� �$�&��T�������o2+�z?��(�K�R�,S�}UY�� ��Ӽkz	�+u�����(4�u��BN�a�A(
��n�{jlo���(X� f�f-W��am9���^��Ne����!�G�>��9K�����\�}�$��nX�w�]Ǣ��v�7\�) �.��$�hW-�n���WZq��՛	�Q?R��'mQ�S$U�����Ɠ��x��-�d���6-��`�����M�+�T�c	��i���ğ?�s2���!�	���5m��L��u�9��u��3d��������Å�A�e���1���[�v�Z�x��ۅ�r,QP�f�� $Yi�z�3D�<�2B�f�A�DS�~-�ޛ��{��"����������%�	Wڣ(Ț|�W�1���V��9e�*��;\1`��ńo������*ۃ����x�%�����K��9���X�?  �+�1Lq7��)�M��QM��!O9�
;�Z�6��ֱ����������oW���>sQ�oՠ�bo���������|��h�2S��-���f�k,
d��:��IoT��Yp�Nw�˻-���[;�DRe\my�b�_��[}j�m�&SM
�NT!�<^�u�::�i���t�'�G����2v��2XG����X�$'���ڞ,��
G�c5_��렱���Qͮ��.Z�xR-��8�OA��:Lb�\.�k
���3���
�Q���^g���69�)fۉ�t��q���+�{/{�-$��T�������3�]��܏�*s���x��᱅�"$̕2�c9�Tm�v�Z��⭲�*d�(Z�� 'n="^r�jrcܦA���s=�n�u߰��7�*�)���S�rĬ�n�(%����{tU�u 鏀�h�̷J�Z[Gמ�A�Tf�\G}��Ӿ�]�U+�~��#$�!Q\�n)����6�|ܥ>L	 mrS��v��n���F^3jy���:�~� =�
4�,�-��B���K^��Z"�b$���ǡM��;Df�$O+�Sz������m���{��ֶ��,���(�Nۭ0_��
��25O���Pu�g*�4ƾM���2�N��ޜ �Q���#��t������ue7U��Z�������C����a��mMN5�i��Z՝! ���Y�^1�9��%�jor��C �\��h�̅��t����9�[���^ch���XK�d4o#vV7�wV�0��C�C�F)��L7�):��cS�� �'UB��^yM�Iё������^&OR�i��*�|�~O���9�U`�ŏ��%6+�e��3����iGl?,�!����׹�1=Q��q���6DT<������ָ����ʇw���a��Pmj��1�/ˮb-���w�M���\ ��	�K	Y
� �=�}��?��%L�85�T�ES�'�a�FlM�j��vC�^+o#h��8#OJ������jL�q�vQѭ�.^�ɶ'��~�����),(� �3��L#i�X���. ��Y�����p(>�*�^�6n���v�.jh-r�@�
���2��v���3@�39U��x `zfA�qrCnڞ:	<�%�����|j5��Rf�ԭ�fw�,��2a%�̖@UM[j-���B�ě��Zn��<��&���Q�=ھG����?b��B�#֥��0�!/�ۧV>C�l,�k	Fƶ�.+ˤR��H,���/�c�M�Xݹe�yґ�vF�I��F
�Z����G���~���\����`��8Mt��cz��k�ˏ�����U�*�e{	|�K*b�iF{�)�����
�W&�qn�qy�R�5��xi/I�ѐD��H�E@8���C�n`���A� �Co]�4�._w�@Ő2\�Ur"��!���cpf:�/��(���	��X�kZ�+��^=6ؗ��Yb�	Κ�ܰE`z���l�A�f^�����egp��T��,:"w��B���wL��ië�C z7�i�ĔG7,�Hm�1����ʥ��^8����6���LZo�����ތ����8w�yrr�*��L�CN��Ny��7O>w��h��)/��a���쒼�3v\_
�Θ��5N����"�Q��H+��G��Ǖ��D�jtk��!~�Q���������ܢ{�u���3 9���㬜|x���f���~�KY㼀�P����`��F&�4�L�s�� ʽt{�{���Y�*��gXN>��bh��	��T�ɮ���|�2�v-��R�6\������b	x��~�.Ex?�l���R�9��1N���bN�mQC�����2��ˢ"j�P�6��!�.�6������`��t`����>�+�Ǳ��+/>
#W�(���/� o�_i����LI�]P������K$�j���$��,@��,f-k�Dȉ!�P3&ұhh���H�I��19�թ 9-I�'`��n��vW��]��XL�H�-9]�o��K}��L���O8 6��(���!@�Y�Ѥ�����X:o��8A��^�ϙ���ZIru�2vE�C�C��3�K5��p���ZI���L��σ��̃�XP������3l�+��B�D�0�7ꞷ�P�=���P�k�D q�c��Uc���J���S^C�#:M}zӾ3��OJ!���+�e{����,zn$�0c�ov��:�����@d��tP�+�*m���flwu�oM�ռ��J>�5��}���@S����4�->N�؆�iC��48bX(_� @m��e�Y�tl��O7L˴�o*L�5�|V\4���Q�-7e�7n��L�#`4j�y��V�uS�@�n.R[�3��{"�b)�%,`��%;�<G�@_�3�3�,_��H](MF�"m�}��F����A�0p?{{o&��P����<������hXH�o��;:��k����x\z���5+	kq��p{��p���:��:�a@���T�;��q%���f�T����0�1�����\������պ2�q���6nD+�����Ac1S��'+�I������0I�x�t�Ζ��,U�<�%2�نrެ���M��#�9a`ú%��9����Z���k�V��� �M�Pܩ[�������Wn����d�g�iC�����2�Q� ���t�3'�]e�Th�qOP#M�ʞ�ք�[/��7W2f����&��B�{�����{����s9@Z� �_y0�s ���]�N1�w��H��W�ZA�{Q�V��м}�������Ef�R[��+8�����r��C_U���#*���MpzMn8^e<��cؤ~���B�`�q��U���E�za�]-�$Q@j��j�8P��Pd�`����:�|h��e�dI� ���4)���������qݯ�崳��'F���4�L�'D<��x�8�9|]8��m���m�Z�yux�
x�/���|9�ƆM�����l�	�}>ԭ?�Ա��&-���]��@�U�����9�qxqcW�+~�ܵ�T a%�ˁ��<I할�,�}۫���^�Zk����o��6)�c��o>b*B�~_f�s�}'�������-���d�B�J�"6���L5k��G�l(J1uj�籯��/!�
��wk�ʐ��(��
��M2�+wWC��/&_PŮF�-�dnLƌ��&0���(j�eN����vs��2�4a���v�y�KD��^�k\Xe��\�6t0m����:�
3V��� �H˫�OyĤ�wMٌ�T.E�ө��C�/ ��ey�!�d���1��,kǶ�S�h*6��1l�jXS�U�G��7^5t��u��@�(�HXE*y�(�{R�(�]gFW�.��m���5��-�� �/ԅ�1�֠X.=�Y��9Lt�Td�6z9��c�1Du\TH�2fI�bSߑ�G?�;J\sHA7�����Kn$��܆�]�lY�j�� ��閪�RدE��l|��3������Q�@׿&$�\���9K�|(� �E�(eD��ݬ���!�.��#�<��A����SG��$���S��2[�>&ٜ ���,9*)m������'ô�G,�QM��P�w�8*�$}*���Q�1¯F�xV/Œ󜩰�"0��<v��7h��P�Q���%)V���M�a��蘼
Z�yp0пt<�R���!����{�2��%��	�E��ܫ���!N���;��	'��E�nΞ|�җ$���D���]+����3�;Dh���'K�b�� oI�3��rt���'~�=��	r�&�?Ӽxm|d!0��B�ה���[*	r�ܹhK����z\ʊ�<�sEy�N�L�<��#���q��Y�|��!�|�'N�s����J7�����S�)��U:���d;��@�,eI�FQ|��Y:�+7��_�̀��%���-VH�K�J׻�|袁]�*�y d���w	��=��vQ���Ƽi�zm���/���:���g-�i�Y��d�BK�0��%�)1?&N��#m�L2��e[������c��UbGH�v����,�,�:���:F|lO��bg��Zy���"����ӷ@����0H�G�0��}�H�}~$��(!W�V��`@�:"!�hp��W�:�Ɗ+�� ^*��7c��Y��^����i5�^<ǄOz?��=~qrtq�d�hw�5�����..���3X�a4�{����q,�n�>�*�I��I��d6G�*n��oU�L/�h�$l���`M�߹�u2AgtS�Wjư�I��¶c��חq<�P1g�򒣜�J����$�.SW���G�E2�6�W�y@�)r��lN]	�?�6<G�V��G{���<���Q�D����������5�f�Q9L�C1�A�g�ޖ�EU�=O���g%�ӔL�&� ,�g�ļ4�y�	��?g�eЮ=�D�h"V�S�tZNK���m%gL�Ow��t~��P�J?����y�c+���T���x��8�)��*#.J0��/�{��7�ĉ�NQ�e*D�I!��6/�_4��qi�����LZ�m�=���q���>���SD��7 �;�(/�'��vrOF��a &hV�G��4����*�3�����S7�(lGI����$��)�� ��S=ѻ���w�3ǁ]�RS=S�eTJd�e�aӂ�I&`P`�&uJT�Lԙ��fJՄ��K|�+<��	̉�n|鯴U*ә����!� 7��f�f�n�!ORZ7ô�گ9n1��t(����]k���=^����#�0O�4�~A��z�NLXu誯lj���XM���Y��I��3��c\)?cw�%>���5B<
����>�G���ɠ��}�tg�ȉ��ڻ�1�P�Æ-��éli�ݭ�¦�y���rq�&���I���NB�)�8�}xr�`�[���4��"�RYG�g�����d��svJj�քt�o� �� ���t��G:�0�K �G�Tz8ia����W��G�V��]��yv1pba�)����K���g���+�Mg-8���Jd��T3&�D�0Ҫ�xC�t�u'c�M��,X�Ϝ����Z}�48�V����L�H}/*F�_��<6�v�a�s�Ug p�)�Z��3@2/�ƫ��n���Ё�3���y�O��As8�yi@ߢ�~�o_L3]ʧ�Zj/��Z��γ1���if���_0ã��n#�� :�ĤF/�����}���M�&�C۴�-�j�'����ch�4X�Eљ�hê<��;�y�h��s*b����i�)�~P��9�汍�[<���qNT���Ӱ��o�-�^���ea���8��ޖ�2c<�D^Ba��f��M&�<G�n0�A������Z��l��a���:8���������j��z������z��)�JW0�5�mGC2�2�-�V'��_�D����s
��2��~?(� ;dY�J�[!��>{Z,�B���$q�@�PR�4�?�15J[ ��ƫh9>J�60e�&�;�N�u�9�Mm���E-����h-��իY@�7�x�\lA	�$G5��'K��/��>����+ן`�6�KX=+�為{܊�_tg�{�2�f1 CZ��:�o�i�6��g�$Ug"M�.��1�������?���gs\��8��L_��߮���%�lCUnn(�������ʆ�;oZL��.�Z�]�|�lBn�&��6pv�>�r��5��B)_�2_ ���%/�Nk�CP֢_c��)��`H��+3Ϸ/�,��zX�FA�V�4!K��_�~B�� p�А��|��X�Q*��Tz}�ۿ߻D;!�A]}=jzS��>��8����	�y��W�4gL�ۊZ���l��C�̎�y�=3@P���������܄XlxV16EB    fa00     bd0A����L��c�������/"�"r�͹B%+Տ��[?��蓚W+�f,�Gv����D�3�/m0rk���6�t��l�5P��AW<N;e9���Y7�!����t�T�-�NC.ȅ$�s��T)^����aS�;fDr�]�{���H�`g#�1Yk�����g��r۳m>�Vh��[�L�p�T�V�9Qa|��S���E�ra��+.����c��7���D6�]J<�_6�B[���Y�i`k姘��ɍ�喓���*Y]����lt����h�b�PiXc����zt�e�L�s���Q�ͻ�������8������&���[�wA!@��²��Yj��H�˝sv��a�q#��q��1u�bªG�����0�SDV��������=�8i�� �߈W0�"�˖���yîq�Kq\1 I�ӛ��PT�9k��Fi�]��T�L:h\�L!qL[�����P�!�B�c\�<�����B�W<�����,|w��y�����5����g=�ez�;}t?����l�Р��6���B�Ō�_ٵ=�����]ؓI't��ߒ�.d�%o��f;�T�z$m��T^���~��ա�;4��Ē,�R��8�(�#;dn�
$�K&3��`�d���@ߌ(��� +-~���7���2��z�3�!łM�Q#��:��]O����$��Ss�&'�bʎ�G��L)���g��ۅ=�l刵�>sus��s�+�������Ü�!�ڵ��<-.>�����	V(W��pdcJ`�M�.]v��<�������P�`(�^$
N�00J1�Z?��hC�������3��c|G��wv���b��Ay��ȼ��{�y��J�U��A"�P��e���#/�R�1�ۦ�b�~�	�{N�}U!����M��R�-�0kϨE&&R��-�|�_�Dqf:kڽ$�r���� Y@��Eb�����x+�����7�<6RFZ������ek�Lb ��R��>��h�j��^�H"<�S���:��	_	w��=����A02�N��=.�E1:�d�P���J��pF9���{S�E6�oNV3MPH�f������_��=iy����x�=�1���8Y��HCm6Άs��]���S}�� �3Y_�A������'�E�)��=�FK�p��LL9E��:��>Kmѵ&���������'"�$-&Y%4���_.@����QrՁb#�o�z!��e(�+ �>G�9_t�	dUfK0Q��R_2�����>��V��f��ަ|s"Iճq���F~�qӭH�G~^�-8�;��̵����$��cރ�'�e7��@��g��"�sH�)��vBo�¿��Yj:��$y����U�2�	�^��D��l����y�ë���KU���S��j����z�>r��bɵ9�ěݪ��ǚD{����l9�r@�
�v���B��l_n�+N�Q�B5�U1Κ��)�yv��A{�B��攭�T��#����1��ȡ��������A�ڏpNV����B徉�Pv�¡9�+8A�a�O�<����n�����>��O�I���7�$�D���=z$��b�UcoA>��%�F"���lI�W��[.�x/ey��a��'�9�S�h�f�����ח'MfW+ˮ�X��R;�����q������>b/d��Ԯ�ߙ�������?�!���G��+�U��{��y����<�!�k���@m��'?i��`�yAi-y���e)M��\�nJ��9j�ax�|��cH^���i&�������f��e�C+ʗչ��+T�E9^D^�>Ӟ��Dr�;
�Y��vS���w����-��W� ����fD��h�Rm�[ '|ڌ�!Z~��@�#͆|..���W/�0g����3��.�̽�]�V�)��`��k���qJ���U^��#�(ơ�L�%N����.�� �P&�5S��Qg,������<e)J�"��D_�/C����O�-D�Iy�@�q�Y6���nЯ�����b�I�u�\��/�Z
ĥ�� 
0>+�u_���z�5^"�O�L^���O�xڣ����aK ����8�;�/@��5hb���D���Iݤ��Y족�,(��u���OZ���km "#�r�S�.����~}�[�c�뿝�R�N�5D��A�'�hjK�+�MlBI�^ݥ��q���kQ�K�zW���*�ѽ'I�t xGVg�I=��y_�N�ԑ/H��C��1v��:ZTø�ڌ���� '
R3F���UFx�We��\���Ƶ��P���:@%���bבQ"�#��R|�\ۈ�V�廬.{-��h]~~H��,�/�3��H}����(]U�����u,���C\�>�cw����R���I\Yw���'����=��4���E}���(W��=%���h�6h��W1���gmj�'���y�z4�`�|��PN���������Et�4b����<F>��hG��[Bn=���������B��ɜ^GWї�ꉻ����]�X�� a�*}�	���#��N��|~����9�o��2��J��x2�Q���oR�1���������ʕ�`7�qc4dev*�����s����[�rȒJ@�J�0V m-�e�,-_�|7<m��F�b@P��I�O-۲2s��I���*q}���}-@M��2��̧_�	v*�o���^m�<����6o0K�ሇ2����c�6W��%��!4H��_�#�rI�/����Dk<��w����(�ώ3�hC��|	#qL0��Ŵ�O�����Y��ɸ��'ab��B&![��&<roK�C<��y����Q�%~#Fdԛn|�>�*�Hl<��8�*;OyX\ kF�"ܗ*��%�a�z�@p���T$��ҫ.�h:y2��u���)��!�)Up�^�|⸄alSmt�-���AS�	�x��=�핍�$�Y��SqlN�̞�Jx�ST/<E\q}����XlxV16EB    fa00    1220�x��y�����$�K��6�*��l;}nU=k_�Bf�޳zh�q�e��*t���#�hr�Oi͒�Q����YN�m��0�(���(ַ��=�E�I�.�u�!&9p\�P,�t���K�D���I�]PPnp蝩z��9#��,/��_n��� Z^6�*K�>!4�x�䉷�»����T��_0�,�Ι�ȕ;�7���!�r�d�j1bzȟ9���c^��J:we���Fn�(ٙ�qF�B*�L�藫��.�����2(@��dK7#Tp�Xv��v�$�pt�{Q��|�{A���Cv���p�aX*9��X1!$��*�t"w�"�Q'��5?4j�(�/���z� �4�tJ�ЛM>����uC����0�9���[a�g������2���!��Vq���d]���E�eQ�"%/��ۘa(�U)�|��߽^��g�:�����'�qM�+�����1�����N7�H;�@���]>�J~ۗe����s���eU�_�� �N�aM��#���%��D 1�|=�S��ujK�v*	>z��nx�ȇ�-�&���9)6�=����=h�{& ǣ��K`��3�̢��!�X�~dO'Z�I~W��ͻ�6��1��>���D�I_������q�{���&�Q}�0
���Z�ZUsߋ �W��;���k�j��0��"��/���m�VFӜ5���ƀ�4��_>���NW ꌻ�$����ْ8�����+��ͳ�:���lP2bg�rEH����=
؀��+��	k���:Z_�N�yZ }-�*}�Ԁ!��u���ɫm�*��D�.IFa���_������
F�(���Su2�3��Yb���B��e��{ApU��������aS��tz�P򒝋��#�24g:ݵ��=��kq9V���!>{~�KGb@��-�}na�@[�`�٥ٓ��Y>7�I4�B��1�m�I���3u��-DIؤyj!�p��<�	�d�<����|Fnh���^8{�!(��O��D�;@���W���1޳ͯs0tT���RS�-%%vp��_� ��F{�:�D$�'�2]��+}�
���3K��s$T��kض`���6��fw�I3x�t2�I�8l��|17huZ�7�\��7Nm�J��-�n7jH��e�FfO�Q�܆TX��>�5�iϞ�ȑ��1�#���wz������ë;ƈ�r�~V��ނ`"�I邈mo���r���3_�u��!9��9�mӱ.xw��l������a��\@����7Up8ds����l(* =cqP�oׅ��%bg���9�rM�a���(������=�c]I�)�#.��_@Wf60G���p�����c�H�Ȗ{\����,'�����p~Y--�ڂ-�v�i$��$��鋆���xX�w���\����S*��saq8uE�4�-iw�P���%��D� Bg�tiw�p['�ƿ�v��U�{K~U8��$�ҀA���9F5��+pB�SY�*@v8�� ��62�z�5͔Z�� $���S��C�3�Nw����N�`}� �HE0 9n���Ex�_�:C��b܄W2������e�y�W�bv
A�aXnD�o/�ݐ��/{�o�c� 𑯘X%��7�b��UWx���SV��S�`4Č��x���p���&���&����(�L>�J�ጴ�=&��\��*��-/�*+�xv��b������'N�TY�,	�)�*D�51%�8�%�eđ����"�	�T���l���o�ߑX�C:�kA��:qL�CӃ@h�Y��5y�)ee�����	�?��ޫ��p���<�N�g��ϥ�`��K~��Û5�HqLǿ*�> ����B�ڑS��ڞ_���(�n9X��h!����5C3��-Hې����Jz��qy0��PI�u6 K����H�h��$E������=����Om���<���7a�}}�p�����cm��MF�K$A�^�fN��¯���0o1`�OB�/%�,�ءW'�܍��hic�Ld�T�Sʊ�6�G�y�����ѥ �Fةz�;o�ysj��sy��M\�O�
��A^�2��f?��d~�`Qz�hcy*���!X͞/
�&�*�w��s��G7�����7�G�Þ���g:��ǹ�Kܴ� 0_�����-��	���8w������٪�X>��dɝ
��C�$_����3X�^�N�'�1L�����~`Pg�ڬ�]�G��\pP�1� �N�ca!N��<�|�[�|II�6GC�y�]Ϋ�o�./�z���#��❛]h�f��Z��,R�� b|��HΔ�@D1e� �v|��.ҿ�
�������:��{΀UZk��w���l�|�����S�5jA�f����ؖ�����`�rI�n^��z���X� o4��5�����������J�xO�`�3�J�H��a��^��������⸓��X���OÏ'�m��`��2b5��%A�#��)��t�/���bg99��n�X���#��0�_ o�eY��������_���1�'K�j�&�v����VǕ�Wʯ�	:��]���Ua+�#%�vR�[�4;<��J��\�]�Q��� ��k��+�.�	�tJ
ຣ��0Έ ��
Kw�9��׋
@k'�����r�����\�� �*����D�
�P���T�n��tE* ����f�`�A�^8`��|ɥ)yR
Fq5#��Y��ǁ�� F�vO]�{�3%z��)���֨�!�ߘ@p�ꅮ���da�yu��8t��灒��0o@G��о��9��S��@�/M�)rî��h��H´VL�1mZlP��4Im>[bQ���#7b=/i�����h�o�8��?�4s�����LFpK�׽W]�Ab�d|�1�_�a6�F�'�T3H:4�/��_��̺@����Ś�!��/p@�0n_Hk'⎄��H Ū~+#|�bB<TE�ꌍSK��@p��.�8�
i���q��LCe�x���F٣s�����#�n��X�%@���i�o�P�HP?���!�1���r��_�ր G'�[]�3��]AP���*�y���!�~_����;��'�Cn��R�N�N|�x��-_A��p��M�ǝ��̜�"�a�p,g��@F	ۿl_~06I�Q��7�^�����ME�������&
54�z��<?�@RQR����1W�,��ީ�:`�D����c�:^���	�=�G!��q̟˔7١�3&�,���2C.E�h���B³�~��Mٰ��F��������y�N{�T�"�jH�p5
����Q&, p�X�l��z/�
�W7j���ƻ1���
.���d�u��^��@P���ƵIE�f^#UŦ�(�0�şT��3�v��T.�$�3s�z[�$5'�`�?��3��.��gXӭ�X�0���<�M�s��:��"�XARhP)QG��UJ��ׁ��a��E�͚-w�����ѮA��ջc��Y�(��+�ԃw�u�;�I���b��v�X#L���o�c����z=_��㟧���m�ٍ>g7L��+M z4n��-����q6���4�:` u l4�L�Az:}+�T:�mו�(*!6�wQ�S8�R���PUM�Y�\.E2�����F��c|Rf.�̏�<1�]:%��j��ڐ�fs�9J���(��W�)�lռ��sCX�2n���+&����i� XL�#lֲ�%��ċ�g�Cg�ɞ�#���B����(�{�Cd`V2��&f)�I���#�j�KZ]j�F�v�ȫ	�$��`<~	q[m�-�0v�[�(��(ܻ�q8Gf{9u���ląii-�݅Gq�$׉�h���qbS�|�	+Į�����8��~F�{^��}L+ʾ��WsZ���N�_�_z�������J}%���.��,v0$���l_Vl.\;-T&i٣�2<5?o|�������R�o	��ݶ�����K��&�+I��hB�����،��Qa��s#�]��G��ź�[L�DO�^� ��V9杳B�����L�P|WD�E++T�2��Q��6�#�b���O��de�#u���*9�K�#w��LHM����$��a.6�L����������A[ܿ��-&'�XlkŨ?J��,�!��([E�{R/�a���� ��(ɚOQ<W$.�� �����չQ�/@��j����5Y���z����؅�{+<]O1-���`Wn�x��f9|4X&"ܮ�!�:r]i����s�O�br�-^��ߺ�9M43`>(�}V̮��¹��:+N@���zH �]�2ڞ��l0�)eES��aT�jW􅦺˔�G#j@�!I+I����n����i�m+m<Һ���x��yf(�2-D��k�4v]:� ��=�z�8m5{��ʶ>!�u'�"�M� }s}�]���PN��d#-�Jt��s'
Q̴��5t3��
�0����ӄқ�J]�)m����C+�H��꼟c��eW�L�?�='�w��n����b=�U��p�v����ĵ7� o�����mN޸C,1ic\��b^�72	�oXlxV16EB    3fa0     610�M����쫰ϕ��'�����)]Ge�L���SDl�X�x�TyE������v><.**ܜw��ou�l'�����5��Πrz_~��O��2۝3z|O����t�99?U�8�qa���y�-�(+vw��%Q.ӽ�x����Iw�m�Q-�v�	�6�!�,pՠl�l��G	�`|���/���=/y����dC<�Q�q�%�������nK��4e��EB��߆�g�`�e�A�x������E��M��y����.{�
���x����mS�pXàưm[�Z�tЄ����r:�EH��Ȕ���4�V+d,~z,�"d߆�)*#��⯯�SUd��@��<OU��"i�g�Ȅċ���Q�L�k>ЋJa��Л�)3�k�[aM9#�c�<k^,��������0KKjȬS��!-X5�aRl���qlgO;Y��?�wt�*9�Q�����__of� Y��ؾv.<��8�3^]�B�h��^����ސ����*@1!NJ�# �D�xP_�<D�0>���EL/6I{VRlc{i.X���!��Ć��9oOk��w�UY�B�$��b���m�@�T�w[$HT��{�Y�qz��JN&Q��%��3uN���`�TG����8�;>��G�\a�H��Q���H�[�z���Y�9�?�#��#NJ���~C,�D)T2^�����|ڜ*b�C���Zb��ұ׋��p�q{��g�ZV�O����{�Pa�2w�I]�&JKoA�q&a��E�����h��TM'�U��p����<�N ��C�������K��y\h��A8`=p���X���<G(^]�E1Ե�[�l�Na	DNp�U+�Ƒ5�-�˄��@+s!�-2=p�x��3� 5���&��}�*kˢ����:�X��&N�� j��^oo�᷹B�t�| �66S0l��3�����SS� ��U���^:��S2SUlD������ߢ&�")Q~�
�������Je/���G�S�
�d$J�0RЬe�.�H����� ��7��E�\a����T�z�j� |�6(l��2�ye9?ټ~G�����/(3OzKF��)�0魓�Z؈�=��{��?n���\�_��p��� ���8�âฦl(��^��c�̵t���6[�I�)F�"�]��`�!<O��쿾5_����bʋ~�Wk�4ߪ����L�A}��
\ϣ/�������⹼~�Zdj�D��q$��/��ۨ��%?v�x���[��ս^�c���uC@���А\N�׌�b[���@�(��8}^+yԀp<؅+���m����!��n�x�/
����%3�	7g!�bBbj��%���W��~��_+�*��ů��O\�:lX[����_qy/�`�m����\K󦘴zSF����H$F"���	j�ܖf�3}������zȥP�X�Xx��yˈ���^ iЯ��S�(*�_r�V��o9������o�a�%��I2Ѽ|,�P�4~�/Y�׫ǭ��ͷ4bHx�$땂������N4
XlxV16EB    fa00    15e0F��@�Z&j�Hn�'{�<;]���5qU����ߢ���Xт���cp��N��R�bL-�M�b�^�2���l������>�v7uѳݴ�iS|�o�u�ܽ�/��_�=�G*8��F�҃ �Y̞ �	�$~#��D���U�߬�&k�1���6+6Ka�������+������'B�U2��t0ɭ�Wa�N�f�${�u5:�o�]-��H&w5x)y�EkNv�\�w�����J%,��ћ�6����I�tw�vD�/��&)`2�+BP�<����R��\/��Ύ�4��g�x��ttv	M]�2a�>fu�K됸'1a����9��\n�;�-Q�#*?.�'Rь��ǉ�.�K$n߄�9d!�3%��Çe� ��z�T�[^J	p��I8�RP�fH0����K8`���%b?w��0�>�9vj�W
f�>3�5��N6x{���	;�R�d�������]�,_�,��?�e������p�T�-)4GW�_��}X����Rk�@�� �m�&5}y��q�]R���I�0��!ڬ�2y�����i���5Q���9��U������#%�e�&��=��'o�h��λO�g4!Z8���e�wU'"!V�
E��wx�����-�>�`*LN 7�ѓa�a�v����g�p�S~[ل�b��+<�A���|?�X1������N��O�/��s]`���!h0�(��7L������j\*s?���?�w��۾3Z|����H:�i1w���9^���NY�t}6��R��K��M(�j�qK"��x����w^�� ��;�Zۅ��1���|�|�M��u)0d}����<J�f]�g>���'���$noq\�1��]~(�'�K�MWr���^��H�
̛(�������)km~|(�x"is)̊k�c��Vl�w��[2uCm�����:��$ �,�[3��[
e�	.�4s���Jb���A��!P����!�Y��:�H�]�%�P������1p�qɶ��9'���Z��۪�bh	�V�����7i��o�B)=��ͅ�r�
���G*�E����o�+k'%�Ȍ.j~�.���Q�5��F�L�+Hr3w����P�~�����aɁ�	�&#�e`az�nĬW�H%��>��4�	�����&Г֓�2:�۷5�ȹ��,�C͖���ӎ�����tL{��G.��Q��: �Z)�\���Mr�W��7c����H����#_��.uiBee|�� IXȻ���4����(Jt�R�r�բż%�\�@�EFC�+����60�/B+��Xf+
E�3�4�d�������� ��E�C�Q�d!Vz _����Є��7cɚ
�?٫s�kI�y�N�E�>�[<��_�O���*J+ׇ�8G���v] w�1_���S&fW8����LD|^��V�U`�����'�)A��a���T݄���2��y�ڨ�Γ[A�5͈Vb���-B��~{ڜ�M��hrO��|1������F�C�{0�rC$�ѰN�����6N�fUֈ�?�I��q��wS�j��dB���m�VT%kp��y�z�EE����r���X3@�S�	��/��]P��Ȅvϔ���ψ�@J�� �Q3���1{�2���=� �86j���Zp˒��"dV�@�v�$�F7�`�������d*��hAK�$m
ǥ�\���t�8�)ϨFT��:���*F ��'K�x;��E�}��FmG�jRH���W��|]��#I}1_��-5J���]G,�Pjl��5�I�h�Iu9�y�'�Z@�iy$�!�`	?���1���{���Qdp��NG����Y��WtVU��J���*PR�K�����ո���V�#"�ْj��w卭�7&���Ņ��սN��-M����T-�uӶ-� ��;o_�� #|qo�Yv~��^h�,J<���g�_g��S-��j`��Z�>����L|�#f��ǫ���a�X�ǚ�w��:W8�hg��}Y�O�̏�������?��Hc&��#T���{���//8��\P�9��G���E���)�Ya��ZE���i3�8� �+mE�{mE8w1�jqs�. �MJL������4�n�L����� Ĝ>XЍ�*��,
�;td1@����{�?��h�=�dV�v�e;��n������S$�C�R��D�@.�'w|��M�}v�����kbH�(E�Y��u��%��V��2a0PM�\g;+`y��4�m��ۃ���>CT~�h���d��p�1��������%�5��_sݯ,��e0,�ZiE��I�����Qkj��;��땧F�~Z{D#���f�m^�*N��3�^p����������{��ǻ:\�P�_ΰ�I�4i�a��v�ceB�,e�~Y7�O�K�mW6�v�֌ �1�܇j�r�P�^��\�'���Y��P�S�ܕ��C���B�az�L܋�&t�����P0���|�,���<��G)��iC�8D=���|���Z�T�=�遀�g���zZb���I� ��q�2��|�j@p�𿨚��y�o�rz�G�j�׏"6����7����I^�n�2P$y�[*G$��
l�'�q��o�M
=ۋZ藌㻜i&�ϵ�S�J��b�_�+�,p�}*D�_85Ɖ�o�uǂV=��X^@���[e�$k��C9O7�u+{�G�CLb��lz��B����� �����n���7�`D.�&�Ӽ0�t��㍫���׵��dX��m��O�p��7��!ғ�+hYs�N��*�^+�š�͝gQB!��,����|E5v����A+s��@�ii��~5��X���eˬ��Բ9 ��%�"�q�"�$i�X���2�5�ɀ�ia�{�.u/S�.�l���
^^z�l`/�g�nOIz/���a
k�׹���\/v�7H�R��?կ$ڭ� �7�+E'nۻ��M��u]��lh�`#�ҿ�'���ɠ�^�0v)1b!f�u���<T�D}�j�+�3���|9!���Y~� j;�o��G���q��-,6���!p��B�!X����~5r-X,��]/�2N~��R�?f����=�ͫ��{�Eƴ�>�a=4"�ː�z�̕1�i��vߵ@��䙵���pP�h�%>���A���7���e�T�^��J}����0�g��(3���9ѓ��z.q��IW�R�3W��󓗣e�&#�%B��B�ה@�Cކ>W��%��]:�xFA�aj;+cזJ�?@u�%P'���K���	��}�w�D}��� �!
�	(^����Y!��ngBb'���3C�}��*��b�#�V�𹳪��X�>;�2������*�YC
��r�m([�';M�S�c����G~lk�
&S9�0�sŸ#D��GvhPt�t��u��^z#Ds�jOȘ�0�� �������-~|tX�i�9h�4q��q����#86�ڣۥt�c���!���AНx? 	\�#�K���7i=N��^�����˦����M���O�V?K����s��Č�U8���խx�����k�v���L��\pnr�o�|�f)H��$% �-f淋��)��p5���i�r]v��e�]͗7M���ԖT��!	о�:�
��k���͘��"<v���ˠ?؋[?�EjhV6+��I)l8�r�;x['�ݕ�y- M��\6U��/�=�Ǩ�d��V���]��NO�l�uT&K��q�s8�G��%"������Q�-շM9mp5�Uk>��T����r�fm)�Ġ�-T%��X�9V�"26��1 �n	�\��Z2��}�)�$-��4.D��-g��
G$��)�A��v�)����rB��F���DB�7�`\G�"������1W�rV��y�A^R
�3%�N�ƾi��u��������LV ����R�Y�wݩf@ h�(Xn���)�Χ�hB��g��,�gШfo������}��W�f�%�m��vB��eXQ֜?�#~���!�k\�/����l�k��7SW�r��Ʊ���/r�;/��Q�Ɉ�"��7�g��I�]2�YIɲ��� \��=ҏe[ڛEM����	#r�&���0g&��L��HA��B�l��{ڦf��A6N�[�:�so��N�/��^m���(�i[�R�!���
�֓@|'s����S�U�>m����#�=��@���щz+�$W�5��"�儔iOM�|x�N���2�}V���c �;���?G_V�-��q�$�M�\^,V���fB�����Z9��&���@cF��*�iӌ4zC���H�Ƽa�Z+<�-1f2h�o�򻞼�y���w,����W{�;*l��b)�U�p^SG]hk���]J�}��{�N&���P���z����#�����-=���3wQ�񝘏LP���;K�.Xw���SpF�����6��:T��4�ܭ�+�Z��K_C~��4L�e�>��X�:�1T���#�Kk7���M�`} td�p�l��'�췕�z\���ג��E�1����x�:���Vģ��J�/OƮ7꟔2�����ϕW�����V�Đ1��04��0��r��s���Jlv����2
��M��X�Kݫ�"�ђ36�}޶��9���v��(
潐�@8��T�S�k.�F��M�s��o%��c�h�@8�XY�E�>{҅��O����z2I���%���4�M�Ӭ,�YS}�KC.��xA�C`�ό,�S���3�{�5�����W��)�]t>G�-��֩���z�[4��< 3���?�..��������_n�t�Qq��I�Х?? �@h�2P���?\�(��(�]�,i���T�N���8�d"�kV�/��#��R�Jl��T�S�=5|����";C)�r���b��m�簵y��������bfg�̯�ZTQ6sA�獉6w��l���*���FgM	N���K�{���8��/��V%�Pl�L�J��6�����]Y����1$4�!tU"�3��Q�#���P}�G^��Ne���H��rҙ�A:vLm�& �[2Kȯ��yZ����X�Mt�) �9�T-䱯~ܹ�n�<�b�RE����������XԮ,W[��Ew��KViI���)e�������#Q��҇���3T�]���O����T�a�$n.E����x�������6��9�۾�(��ȭ��k�]��hg'ò�(�	�w����l��Q��-x5k�������83j%L[�۴jJP�"�k���*N�˪iE����n���Q]u��oӊj	��3�a�C�1�Ct/�#���7�U@y�&Q�R�!��~�3wF���7�b��$����g�Q�/�}�Cp��-�r�<q�+�'6͠t��ؙ�0g��%I"�����P��#<��,���ۼ�?���n��X2V����t�����c�,�u]�)����/XlxV16EB    fa00    14e0fN2@�$
vb>�l�O}������B�"�&7��HV�3[X���L7>C�ю]mT��͟Gd�Û�m��~����yQ�Y�j�����D�� el�QM����_p�8~���3��#��T�����*M|z!��뺒w�o?��� ٖ:zuL("�\8����g( �~�=��'i�
�?9m����Ak�ye���pG��	*�f����9-����,���Ǎ��\�2H��F����u�r��.�2R.�M�^SP6/8W*�\O�~��OVY�:�H`~�][�Ln�o�T��FJ��g���Ý�u�Y��������Q=	z��ms9��O�f�8������;�o�%������;�G�M,Ӓ.̥�|�щ��TEl=	-�+b���c�f-7wt��(u-FM��'������*|�)E�Iї�Flt�梕�Crk%Pw��s�|,��{o�g����>ȁ��X�[1����G���x���!��[WWA/�ɦ[�#}A	խm�QMMdш�*��4�Nx����V����W�n޻(��j��?!�P�R������� �@�FpI@*
�
�2o ����I�Ty�y��o�ܙ�*�r�p��$;y�*��!�lU�0gPщ�a��W�åeۨL�3����L�k��pI	g�@!�(F��ى�Vo�@io����P�C梺=ַ�Q�{�Y��{k��A�C��u	}{��m�}��ջ�
�uС%������V���z��2ܡg���}6�4�tc�b�?�~�@+�sԷCV���(��lٯ�-^}�<d�Vd�r�����p�.�j��\Y0�W�7� ��f[�\�f~�.�5ڢw(w�d1N�O$k�d"=u47	�=۰�J�Q6�����`��� ��:����l���j� �?2;�<���Zd�[��c�M���C��_B��U�8_�0G�7�٤��藻=*��ȭv� H��Ts�a��D��+���׎
G{�Ht�i��]��4a���3�>d}/��������$�5D�9q����
ܣ�gs�.���3y
ȳ�
=2E>�[ۊ��T~q �|f{�Tኟ�鹠X��& L״�,R��0�s���:�Up�/�K�́0�j6��y��|���9y����EZ����ԑ͊Fm������e���*���zە8Z1V��\}�3ɝ �؉Al@vE���6�9��ZF1�#V�Ȫ7�eR�@>�V��V1�,��l"n��P��ؾ�o���l���2��WB[l,	hyr�tŻwЙ;�K�I������ٛw��ۨ%~�ߢ!u�N���]����pjx���=	Ӹu;�����QcV�?�~b�^ffѕ��@{y]���.�Y $kp�x����˂$��&�QDx���ԧ{z�(�"h2u�����y�A�1���J�h�	���Vc��P��oA�� �X��������u�_�RDI'B������z�#�FFk�dp��/�~��%����44�����*c��D��K���#P(Z�V*:Ku�d`w0��j���ݎ��紙�
,�G�lQُi����Q���,nz4S��[����饑��|��仏bO�Ӥ�FL"Qa�8Dީ�e����]孝X�6뢇"�`��GXYl靓�ߊ��|��}	�����w�D��;_W�,�|H������n�8�P�wV@��̥�u�'�Z����Q�G���c)	Rr��tcq⍍�G� 4����/����0)�=����AY���"
�>14�!�j>I8	�0�k�*�� <��6�iO�1խΤ�Oh}��5�J5�,B�q�3�@;;��s���_��0����6��!����3���}�6Z��M�e�3�.���9��{�<V��s� -*���v���
�Ճ��vf�n<��K��"��"�J�hH]��u��^k�����~%���K����D���F�[�(�D'�0�:�4?!�hq��CY���ġd�� �t�~���`Bz�����N-�s�8����t�8��k�[�L�o~�*�f.on��lk���F�k��0�_w�*�,yg��W��������^?X��b��<i��E�T@��t:$)~���?��1�KG�_r/���I��RW�Gpשɧ%v|H���X&T�Ô'[T�ͷ���_�=�����w���ІQ��f�I@���PҊ�?��]����BZ��W�_����BW
B�F@�!�HUmϯ�N���<�9�ż�>���N�&�Os+��v��8�6�����y���C=>�=m_�)��l��@��.��K�zr ���5��(1���(���ƍ�\�.��'wJ�O���^��Y�mU`>O7w\�x4���*E����o�Չ��/Ct:��PZh)�ɘ�~�_��5��h� ���{�D�R��i���K?Eږi�-���TpDn@lԫI��Vs���f�_[J4'����FmCl��(d�.
������t�l��u��R�V:a���i��PM��L���α%k�X;/�7,V���X�7�>��Xް���P�쌉O�T��4���O�A�����EF�ϳ�U���R]��"�x�?n�i"�~k͚ܠ����%�!v0��Γop�nX��Z���ɍS�4����aGV0�:{�^X�:[C*�ƪ�$g.�:u�;�̭ʌ=I
'ywXկi> ���y�J�9��73p��#@�uEx�?�iY�(�Q�yX,�|%�m�O�������G�_xR6��F����3x�Ɩ���X?Ī������&?�d7V,��G�%��a�����DQ�^>3K�IR���R��i���,�[L«qұ�B8#�"�q��İ��B���R�r��>"� �C��Ѐ���
�<6�6rz={�=:��t��^�7�dK���=͹r���G/r ��Y04)&O�ϮdDǵg����	�G�.��8ʁ{���nTq����^~q�v��sH;����-6Oj�DZ??갊�߽��SV<^i�~"C�<�a�R���}�*bĦ<�1�:�͌5'�D��0u�o_ۍ{��6��2��,:��v��w�7p��`+��,��� ������@bJ�<TI'G�P�a�1���>��t�U�
5�'u��O�K��ٜ�%�vH��,x!fC7�"�u61����@�I��IeZ|;���=��O�&?�K��m��=Fh�����I[��K��=3��]��F}A�cziʳٝ��+����ˌ�&��,}@��LG=1~t]b4qu82���O�"���A9C����.7@u��Ă��4iaoƈ,�=e�f���:B>z��s��:�k��8���/�I�^bf�k�N�x�	�"6TE�>�A��]�4���4�z򕶉;�n��]^�;>n"bJE�>�uBhm�	�tQ�!����[d��[2k��΄q0(.����a��{�N�j-	�4��w�<jT�ҡ6HQt����3�pYb�-8k�ԅUy��*o������s{�ݭ;�Y���l�Yf�D���g�/�����Zm���/�z�}:�e�!iLHS&��%
2ȸ����#�0�5�U���km�Q��і�;����>�����7Q���xC�IY;���b'����N���,��#�ڔ�vLc쵮o�D����������2w����t+�� ҉���,���B�C��b��*�q	�v^�&M,���N���Vԇ?T��(���rM�����v�����Y^�o�3?-�WL��$�`�H���)����ti�oRs4�G��d����m<$�����mN�_��4k��O����<��(o�*ވ��fI����5T��ʵ��ݓ�	Ӊ�����q|-�&���b�o��/G��3F9�����r҅��r�8)�P�:a�YS��:C���2���q��T91���R9�},/B<v�������Xg̳4�&���h�,�Nj���?��-�PcO4W��7�'�i�;}�N��G�-���\�p��h=��x<R�'+��!�VTP�.��f,�X�C��a�n�����|�� �ӧdg��W��ī������o/�_� ��b� �?Aj�,�X�?��i�)�{n����?�2ߊ�8���/�6��C�!Ֆ��[��6=D�}?���EK���4�o�Ɗ]��=�q�B&�%xD�9Hg�g}��{�*rg����y�g�C��^Y��3�
n���7��-u������U�sr&��&��iI_H��&N��ٷ>W��hgMjَ���������6�D��Bfj��87�?��1n@����
y��i��I�����Gx�:哧����2d��";�Npw7��Q��B�#KY���Q�O����.�Բ�>i�$���'�c9�`�B0���&r�fb���=g~��V��0��;�]j��<n$`:r��7g�(��^-*8��;��o�q�b�[(��R���wD�XD��?�<@�Fz�~M`�4_��d�W���I�?�(K J��� v�h���}��wFk
��z���@�}Ғ�T�ҵ�ˊ+��.�ߚ��OC�-iݶ�m��/�K��> 5l�kf��7-�����dx�|�(oJgC�O�6�uљ�bg���ЈJY�5�gLI��ZBm_��f�Nj��+� ��H��߼HS-�y������Y.�����SP�Sd��f 2��#[��N41`Pt��nlR�RiHV��܂1�>=�9[���������<�·(��L��֕�!�6������C�3(u\5I�2�P��#fb���0k\�?l��F_e�NQ�j+�{�'��o|8�8�POսy�]8���y�9��ȱ�U�t�S��M����_MO�r����W�׾��E %��Hm���ll�踓X�x﬇�~�����[�{�`'�ܮ��	k�>o[�qq�l�X���3�'�51!�@,��<5�v��A�Q� ��i��1�������TƧ���?�d-Q��Է���}5@�G���;��&�T�1�O&6��_��ȠH�s�	lL��ks��I���ًY��Y���]t�V��~Zb��w������Y�]�L��Os�]�����'��{4,���6��l���פP@���^�/��*m?()��EG a�b3�x�l�{Dy9����a#D� L��C��r*����l����܍H�x�TY9�M�^^�\���J��2Y�����,���ã�f?�+D\�����:J���hҝ?XlxV16EB    fa00    21e0�a�"9;��EnU�8�z�*�����
2� �����6�.J���9|��!��#� ����N�X`�Dss��O��6*�͢;�^P��P�Bk:lyAY��Z�3a^�Yg�р�Ѽ�FÖ��'��A���6�
z�a�����F�V����c��A�f�A7JW���?���w�����yt��"2߉Ï��"갾����8ĥJb�_���ޏ����".�:����?�*��cj~�%��ﰶ~�K0V��P��;�4m�x�"`���
����<��Y�J����a�34��c��l:�����,�SL��w�ŕ�����H �0�,��T�C��b)f�Q��P�����T�U9b�&��6��l^�����!�*�,`��"�y1�t)͂Ю��r�Vu��ך�q�ݱ!#�2�m�����b�w�%��OdU}Z0�Y�x*��/b�ֹ�g\ϣ�u/>z?'�����ǚ&̎��Qa�=��/�\��~�X��S��m�|fе�M<�B�!1���H����[�A�����j�/��7�ްY����;J����m���lE՚Z��yr��ndLg\وƐ� d�ʫJ������D h1;�&�c�>���;��9�O�QP��Ӵ�ɋ^;8o�m����O��Ɗ��j��AR���/�i:܌�թ�%�L���o���A8`-DT��Yݍ������v��v{w�����{J&JG�ҁ!L�?�T�0q0@$�g��t�Oi��&C����t�µcH]�g:�S��^�8a��n���>�o`�h��G�U�n��S���얇�d�T*�2�Gאѥi��믓]R�����RP�}*�{Ol��5��V��ulY���ͬ$��3�|�&z+��K�����`e�O���PJ�G�p�h��
&����w�!+*���k^��c�|T�dY��5��(��9عP1%�# _�.���_R�'[Qp���L�8�8'�^ڴ\$���<��x���]�;bmQ�YH���Ï�W��h�g���5�+��xt�w)�-��d��8� �s�0�06������Nd���V��GI��z�+�v��h����7���~w�rF/�;����-]�R/e� LSTi���m*��;��i��cv��
�jH�d<,^�7��AQPn�#�Ϟ�}�-�mv�-��;&i����f\�8��`��l�(���r���h5����YE뢩��I�Jk#+�`�U^����]�t�}IB	gl��8�Y�by[](8<�P ��*�G�&4Go=MT5x�
Q��?�KJ�AFZ�t>vL�Ţ�~f��K���H��;�D9�_"�;�쳘W�ǵ��r�R$$S* ��#��EH�����sW�������̶���Gc#�'w��rLF�ؙ��<�#��IgI�4���N�������ד+@p��������S��
�R�
x��~�!I����7Xd\���H��f~a����� �;6���ҋC��|C�i�L@;�6%!�쓑�F��^s�j�㮦����UG�M8G�`.�^�)� ��,��_=��PWɩ�� ��<}��?��0��^���ߩ�դ���1�Wu�}����Uݷ�w���Eh�'���EN$���{��w����Q!Bmg����?�J	�ک���9��X����`9����Y�������!v�����kSk覉:r�����?��	������o�ϓ�R.H�û�k�� �
�}����O����s|B`�O;����V���A;��S]ml��Um��<D��P�$�'?�����X�%�K
�[p ���(��GSX�����;��ߖȏ2�����F�)��~j��8�*OkƓ�^��P.ոg\-ϼ��u����̉HEB\ψ�P�(o߀�<�5H�S�Jfд�:�X������So?�@ˆݣ���.��b���������#M��ԁxP|�l+�H�k�L�ُ��~�T��2ulr�f>ܱy����V���<��� �aJ:}MpS�ĔpX��4ڡh��1�D�5�{��n�i �H���͈\AF&����v�-��D��]�twQ^�����_�E�8)� =��d�M��l�K�&��QvK�-J|^M�Qn�ZF_l� � �F��&�,�諚��<q��	����L��A����3Q*a�Q�(�`V� ��J�޽m]l��Ύ����.Osi����L�ilr:ӐBk�>$������~�g>?��\94�Ћ�>44��9
>�؟WI���&>:��
5���C��"���M�m��>�R�`9��Y��S����n/�ۂ�%�A=�jlaæ�Z/D�����$�#�5c��e&��$����{��5r�lt��gx8�R�Y�u�G���ŏ�C�	d����dp"#B����+��O7<��3�y����y�C w(���4
�k�����<fˌ���O�\9���*gOU� A�RS�2<Pߘr��f\`��k�&���O�'�HUs�`ꌜ*�\O��o��k~���\΍
�9�/��;b��i�n��N����J�����<��}�@S�uOa���C?b���ͦ�k�h�J�,��L_�J�,Z��0_�h���IY{��]\��{,���z���������5�J�]���A�.oe�21��K|�ݐP����u!�&�Fp�=$-��B����C2_�R�&��G�@=G�$���] �tdm���Z�X�P�F.�cJ1¦�Tf��Pu�ۚJI�.s�/Ŵ�}�:c�˾��>�W�����{�9Tи 7��/$���&oP���ܡ��؆-��e Iubm��g#C�o[��-�&����xY��^$v�T�R���y\���a���	�ғpPf%[�����>y��[�r�򃺪Dn�L�f��R�(i<��	���U��8L�f�+[�c�r��:N��ᰶ�d�I�6��%A��|�/!]���L�c� iC7�CG6�r"�K5�����?��@�&�wF�Iv�su��W�z���{�,֞��ڢ�D�9��Hgt�Y������P����rĢ=�v�߭�;�RT�Ot`[�{�_79��K�'ԋ�{�)Zt:�>���0L�N�S�ʘ��]�Or��(~�7/�N�$;�Y���+I�|�������r�bϾ
3~ԫ�״�(Q�[]�@ѩ�LJk��1_�-��		�"I-���iS��Ij�&�/�5^� 1X�V۸]���bv��D�6H���^�k��S&jFY]j9��6|�yu�r
��R�y����>h�u�6��OZ���F��8=\�ٴ�x�ߤf��z�B]�y�S�u-��.Ɛ�w��%��7db�=(Rn��0��H�ep����]��|���t��	��G��lrYG���'�pL�H��C��GP��;S���K�y�,cè	�3�<&dj)NJl��IG�!||}'?l��4ȅj=.�����|�9�ިП��}a�%��
���U"n���z1Ā�X�ڐpo�
4?�ds���J�~(kj
�oJ�F�d��9:��ַ)ǐ�'<�ƝJ�*���ʌ����S8X��������:˭V[�h��:�N���($��!y�/�����T�>yM1WXR���}�-�
�W3��p��i}�|3�Lz�'�Tx<�Y�!5�5Rt� ;pUuI��?�G�=b=3�:�vp`ZU�J���Q�$�J���|�F}F�klȣ�e��rĲ.}Ǝ��.���v8���p�V��:�"�m����f��:�|2�ʕ��#��joS.l��:�!"m ���E3�ib�^p�HnL;��n�*K,�V�,	o+��ƶ���"��xH������a�p�`��Y��f7�3�~��q,��2"�/g�n������sĵF�S�d���.6��,D��i�w#W,�g�h���o���a?4n<Bk^5���x��^B��m3�u����1k�Ҋ���p��Z�Јt��a�*k(mt����EVj4��g�"�⡁��I6dӬ?	�Hͬ���-�K�(��k�"w�I������/TL����tB/�O;��`��� �yW��ȷ�0�w�Х��D�MS̳}h]��-T�0!��a�Ӗ����Loy��(g�7�ln_�⽼��pV3x���^�Ly��j"T~d��)���Ҋp����ZB�0��+!�O�����x9?���
�l���|��}�z֥a��
�Y�b�W�,��O+%P�����6]�wQE�C��ܜ�.�����1b&V�Io��|�iT�W�ҏ��D�#�4��Rf�ǈ�qq(؃��Ut��R�ิ<��GR�Y�>�YD�ډ��J�r/7�3m�.OA/+���<�ZAs�A�"ڠ>*�[B��ӧ��.��) r��������Dv�nD���Y�h{�~�W0��8]�h�VTa�;=3���v'���Z�虱ٿ�%�̱�����*�@���[�"a��6�}��u�G�Z_�]�O���.�u�!V���<K����m�KS��ٌ/`X��`c�����Ң�M�|�u0Y�0Q92"eZ��Z,�����U�;'�aT$ب�1�^Yo�����0�Γ���^J޸Y��ͣ)o�������+�+��	2�#;�O�����jD@�<h
�}�CNt+�����4B�.n�M�#��:�J�=��/ҞPq��޽y�9�H��Uќ
���G�	��Ei]�����>���N]_k�-��Ǭ��ZE��Jk��j�gmt�a�6��Ȳԉ��"��Q婩ڬ�z�'�R�%���������"�;����A�)�#w{���:�Gn��Յ)r&�?vI�����k����ܶ�Q�z6��eT/U�~�/��j�!j�}�^P
��;vX�dj*{Pt�*3�_��bS� ����)Wk������˧�2B�Y=ZID7Jp"Z�,`���}{J2�G��0bb�Y����T2f�ai�4O<�����Mr6��;�%1��}P���[~��E��;S�X�8*P�p���>�UxP]y��\0�&w��[�U�9cv�40�U�ڀ+�)X,L��+"�i1d�c1+�?R膆�i�5X�O^����Acp@�p��L�6-"B剙�H�T���3D�{��yDJ�̙X(EL[��o�Տ;�ē������G�|��=t�t���jz,_D�{�db�ň��r��Ӿ�%��������$?m�{��	s�%wp"R.XM�	�$%
��C����6���:�[T�'�z*|x��ļ�F܎�N������o$"�<�S����a�Yx#Tap��p��т�я�
+y�r�ϧս?��04���m #�=`7͛��v�"���/I(Pr��^ 7���
�<8�u�
�w�,	���~"���ᶪub6j<}F�W��u{%N�ZːM9������|^S�<�J^t�����[+d�֜IטÜ�-wR��C�Z�]{�%�b6w(B��a-�0�bgr���s��u��_�o�Chpv�4I�ܫܿ��Q`�P��ݷ�K��K��dTcObf�H�T�y3�	y��ɫ��"�oi(�R���*�r�b\�b^��� <��ޔ��U�I�_L��Y�+�bp��o�9'�lO��e�ܚN�2c6տY8*��N3<W+Ld\�b=|��lz�)�z뀺	q��
_�QߤE�y#��h{�|���س�	!Y�Ssg�	cő���!n�-��	Ew���[�:�����)�h���8TA9�QbN��ь)�`x�:�㦯�\�o[

�K+J�u@�u��c^T$}�q�\R�����DfEg� �;2R�C���2���$fE�]ɺ��6;�:j�0J"��S�K*�������=#��es�D�څO��>|���w�{ĬW�"|S6���t�-3�F)ú2៘ɇ"A�G�V�t\��nnJ!t�@��H��̢L@����+DK�O�����<8ܒ�*��j��Ay"���QjO7�y�(֤�Wl��}��$�����U�s����~���S���[	���Y(\1���Y_-��I����.E&�+�īZ��7��[�Dt �P�DJu�8g=[<��fv�7�|��n/�R2�L�A�n��X8�#2ͣ�U��3�� �O����Tt�@�W��5Guz�����w(Ss����X���T�I�HF��O1OZ���ӎ0�1���q���~�ū0��fy�i�k���@Bɒ�26�"P*ލ��DAw�6�mO
�D[��;{�/�'��X�oo>��q�Z0@M/4�f|p�y�!�/27�+�>�[�y�,=�!��=9 �4�qN������N/j�j��lh�R��B��m
/Hơ�	�B�_f]ڜ�0��s����~����������pNA�&��Zע�>bQ����D1����Ɇc���RF.��r����k^\w�uNG�ȍ��K�o��6@tx9����1�]&��Q������9�Ԅ�P��t���w�������]��U���g
_�U)�uۈ�Y:*�|;:�D�0bT�_��P3h�M:x+l��x3�d�m��5��������? n,��<��Q�k��6�\���I�%�7	:�-���j���~��>�G���2nj�4**���Y�y�Ek�.l�N�ŵ����f���{(^�qR��] ��C� WOY���k��#��U�l�7�~w1��
�L�pU��%;�F`��+���d�s�ȶ�l�l�{�X�|z�PH�k�E�L��5(������OۺQ����T)6��-�d���y W�2�����MZ�5t�.�Օ���ҕk^�N`��^2"AϮ� �l�Jš��$VTV���po���Y1MNO�^C�U��VB�߳{���=�p;��L6l�T�_B�TKOC.��.�p��ռŘ����	ׇ?8w"��T�$W܎��SI��i�~t�-��>�.&�G(c��X� ��*v0��R�[�~?���S���D�,;��e!�^����wHm����M$>�K��V�nG#i�`Rg"n8a�g�	���b��x����bY([K��VZ.������UOz��C���E2�y��5���G���؆	ە3�.>��h-:����ܮ���(.�G#�(�8ub��ک�/K*Kp��˧|b�_iLO��X��`t�~Uy�dF���R��4��n
�v=�t~?��U��	��%��Q���&�-V���b)��KDQ٣��kƧa%��'�[��C^�5����o'�����;ۺ� Pvz�m��L���L�<
��L<ߡ%�����B{p;x@`�gp�\�S˖t�>n4�A�r�dǺ�ܨ -��ﱝ�Wq{P�Q�ʡ��,�n���C� "�Jb#�fڃ���6����pZ�W�)�4��=�HNΒ�'P�����JB����ף�-���9��J�4xT�	�{�RW��s�d���(���h�w��Q������hr�y#;�a{�Ⱦ��6��o�!��+��,l�w��)2��B�mE!�=�ej|�����ޅL��	�i�����;Q˻%E���>����"vM㇒#�s�V��M�r|���MƐ��qw�W��A�X�J)�5c9[�Y�m�a	����zp������@8�#�q�� N�&��=]w7��t�جd��e.�,0�M�ѷmE;�R��s��dú��VJ�C�I}ςM�Lqw����^7�3V�H��Z7X��{:���q��M��(�K����ts~"k���Ec�g�PJ�D�>V��^�Ne��-�>�܋D�I1�q,i35�6z$�%���1ac���P�'��wqvE��m�}�?��/!����j��f��c�sF�^�ƭ]���E�Ԫ�a�N�%x�hu�Y���	��a]n����B�My��Vu�>˙�Elr(ҩ�X�?���+��o��r;(�V�屦�3�H�U'�����9�H�M��/c��,$s��^��TuY6߂�+oǯ�'v32ͫć�O���.��&��N��eRc-�O�L��A��骢��$Ȧ��}˖��KAs/����2�4�4Ń,��c�~�������׎a��L(�I^`�S9��"�6=aQ�SV�́�\R%n�(7��Jh
��Åᡜ$ĳb�a3��:�};>�����A�q��6y\囵��"~�9��� ���9e���{��K=���b�� �}�x�h��~s.h��-(���9Y}"�jtǀ�o� �@C��M�%�]��IeE������Ђ�=��f�T���ưTXe���a��"�N+�
N�i�-<C���!��m+YR���/#�hْ`� �(���q|c"֙璂>htE�O�����2�<i^mќ��}�MkG��59m��1T�t�oOٳ���H�:*�#j�u�gd����e3$9~༔+Ua�����3	���?��B񩌻��#�T��v`�����#Zh��j#�^p������T}��*+Y����2�*������k8�:�P�V�X�r�eA���\x���M�fc+��/XlxV16EB    fa00    2040�x)��8�W3�d)|Tcg��!K��֞�X��z �=0��T���o��X��U�ER ��8�z��x�1�yD�y�:��5��N���F{"y�^*�LZ~]&J2���M�:�V陁�!�L�Fp��CP��eִ����>���[W���	�Ց˿���*�����2ӥ-��Z]&���ǣ�W��&��=8�q~���t=}�v���?����ڴk_zv�mI�2����vϐ�!֔��u�._�)�]뵲g�u��}j=]��#�gP�C�q�3���B�'A����,!��*W�Uླ�A��ވ� k9(���P���tȤ�=A|�	t?@<$c2 "(������II�ņ'[柧�j�2G) w�a��j(WmҔ�X���@w�jS=epiȱ��0�M����}��'����ʑ {�[0�/t��eY�2 5'��~zsi9�7�O5'r���=r!T��텀?8\����T~bӴ���������pa���^�HY������{�$��K@}����['�@@����F�_�'$���rPHOF�;9�;�D�������8'@��54��z9gN�̒4�i��6�aCD�\�[�R�
�1�����)b��q:��Z��x�K8�7eqjvĂ���zH��mUӖ�3�%�6̂�;����:DE�t�d>H���t���XU})ޅ�~H7��=~�i�~e�z���&SEAC��+�#�ꑠ>�7����ߒ`��P(�@{��X<��p���h5s���Ƌ�mb�9�д!��e��SZe�קz�^O�m�\���N�4nBO���s�D���,
�����ä f�JA1+�������|�TMB�)�z���X�������V��8�d[�NC	Rܶ���Q�V/��H��Є���O�(�1�D�U *vB�]'�U�Ú�c�H��S�������m�1�t��m��{^����g�H��SMނM�v2G��Y&֊��!#!��UwJ*�d��Yf��D��ا�z5�476&*���܏[Td��x�G&b�V�t�A�ds�GK�l0$���aw����o�����+'��i�FXξMI�Xu�W/ 2��v��B�g�KK'��(�y��w?�24D|��>@��M��"a�����:��Fߖp�"�X��oU�njN-'|b�ܸ�c��Rt�Jq���|�4�rW/~3���$+P~x�FE?Jt�W5P,t�kx0'��?b���� �iO�]s?$�6WE�����m���|M{?IĲ�Ȍ!���Ѥ��&)�e&�~,���sߺ��������+��$��T�h��E@
ˈ�?a'��3gǫ�j��d�
U$�����	�A���Q�6:��`�0�*�x�2���\j���\�%�\s��l�NL�m$�.����!ٛ�Pg��\�$�����s4g=��w�<�Y��?��k�Ftfo���۔)�< ����}��y�N!�(2WE@&`O��n���P�{Nv��i%�f�������'k�X& _��}��*��>'��S}Ǆ]z����9H
h���Ϧ%$q7dZ���xx�����0[�˛
=���Yix���5׮~4�%A�߲k&�x7�`F�rh�]>ኧ㺔��?�����N7=v
��^2��H%
D���F�F�eq�7�<����̖���6�~�{4y�� �O��%�*�d��ʶ3������@cՍU��;�b"r�`�XzA�0#_Rq �ͬ͒	�;���l�2����(e~F�MgYt�n��Dp+�)��R�7y,��-���=>D6�<X+�t w�b�Uw^�� �q���B��~��˔W>Jݫ�������?=<α��,������1����M1[{�����B�>J�Eiy}��:P[N�D)�367 ��;����]���[���D�����p�][�&�/ݥ�����s�w-<GZ�8bڱD1�<{�0���Êh��`&#R�5.��3ry��^D-IX��/��ͦn���jM�U#�X��e,�q
�Z��Ԧl#b+!H?z�9:�MvC���E�^�lմ���1鈌f��+S<-~X,b�s">��9ONIrX����Ц�`#d����q�S{Gp�v�?aݠ4��b��}�s`}w��2���iڱ��U�ܷjs;���Ϣ��P���|��7�O��%��F�t%����8�(s�Nx:���s�
�z�a?�����q	.�զ�[�?kĉq���{I�2G��}��~�_�Oh��"p��ͩ��
v�yimڝ�R��\����~���W��:&�X�� ���`�\��9F�A�B̆d��_Q�}��EG屲�P�6Y5N�6Ȍ�~5���v��H�`��N�B����ͥ����m�����F^I��
Y�c�7а2�n�|��qG(P��<�)e�IK[]=�s�$�q9��J�Ƹ�[�hu�M����w�M�����,���D�����P�e̦�Ǧj�����0v8�0_hk�F�k�#D�9ΪXѪ��V=��������.3� 0`%� HL��'�*H5;�(����"���}�$+�O?�9n?���`��e���)����g�����Q[�����1]!�|�ɤ�%�I~����x�ݳ ��@˴�lYi}�����CT�t��#��<�w&�����[)�� z��Wr�I���y���c &P[���.=��S�>�����{�S�����f�����j5*s�D4�҉��w��b���>��dx�K}�j�Y�29,�['%��<�7z�?��6M��~?��I����!f�k���/L���+��x�N�=���2�n�:j�n-�L����07K^E�lW�����^a'�����{�m5���]�ُ�䔞�j���)�-���^\�M�9�w�g^7y(��e(I���X����3nn�m�ҹn�ϰ���sr�%��#A�,+u���0�QP�+<�ݗ'1��"���KO��_���m�|�&��"	4	|'�龊���Y<�7]a�8���T�"�YoR���R� i6�^�!��R�k���j�*�.کyD
|�{"��,��VG��J���ӻ�����lZ�m�C�]UŧS$�b4=����c�VT~M��;<l���v�K,R�
�9QQ�Ɗɬ�xx����=b��B���h+G����t���\��v��lq1���B+�Yl �'��+��fU�d�G�?4aKxKvf���30�q�K(B�t3#����u�r(����l\"^+��󢩈5(약j�?˙=i*�?���V�Y�Ʈ"��g���ɷ`:����˲<xW�BE�A���D�5�w�o���1����җ��R�%�N��ط��)4OB��D� ��_P��.�%c�>,S�H��&�d׆��*�
$��ql_��N��O<�i���Tm�E�pwu���.5�L>>f��I?���⤌�"Mēw,*E���1�|2�X:_�J7��b�d�yc�ǕU�s�N���� �~����t���� e��Sy��߾$c�E��W�+(^�V�������!��t��̝�X�H�M��Ρe��7��K�w�'Q�V�E���.�3��l���D(Q�^�x�s!����!ϩ&����g
Л�G��@}�}>�K�0�,b) ,��g��(�5!�B�KV ���'�L,.y{��?5�=d�
��iP�~K���Ƃ�`��KZ���#��{|6{��y��V]�60���~�eQT�/��, =�I�f)��Xgj�Ug�njSLFCi{�[.9��p���r>�_���q�D�5�v~�Ύ�!�l�Z���i��ާ�s��,�<�Ou?KD����6Ji�N̨\��8���lx�b ���NФI50�Pɤ�_��H~�h����(�R�{c�^���Py�Лz����쎂�Ǚ���8/�+�@�=�j{j�w��"&��@H�X����e���Y�x�c٫�k'3�B]��$������V���f��O�ۀ:NKk�eI%dr:ɒ�=Q�G����`�j�4��X�+�q��"�����x}�P8���*�X'���h�v��yFHf���rc�;yk'AY�R�I�Q��d�H�M�עZX[�/�����_��o�F�M��c����|�<�׺[�Ov�+?ge�v�4t#�?�=��v4C��5�j��\^J��?�����<���������A޽���v	RoFd�yjf�w5 �Y��	�ӗm7�n�"���@�#u駚=!PzP�E�֪�4��37[FG��,N:2hV�6O9]i���!�T�8���DE*d&Pu`��-T l޺��PW'(�n�V���TtW�qe�N0�\Jġ� #�z�q'yj^	��ߖ���h~v��Ć��7���qBt�Ts2��U���%E�L�йGa��3�@�^/�H �;蕮���bfΡZ�=��Z+2��{�s^�S�Li?�Df4A�)�K%��0L`b���6�n�"Ȫ�I���>"ر�����?ќ`�*F��z=5�Y�}H��31op�r�;�Z�Kt��k;��Қ,0v@��A1�V;ļ�l��ҹE}D����l����B	?�]��ȧ������j��j�R�X2>B둰����uJڪ~6� �L}m�]�E�L�8�+�L������	�6�/���2�'4���kG�ܐ�����r���5��1%��[l��K~Rs[ P©&1Rf;��q��s6ZZ�ܪ��@2��>:�h����(��[v����/8_u�#3��GsIZR�Qw���d8D���G�D���2��T��|����b�>�e����o#k���x8`Lg�T�	.bX0S����<3G[��L乗m~�o\s@J4��`���F��F�QL���5w;�YD^w﬙�-���=��Y��^r�n)��"�}Q�G��*�7��:3�;�:j�cm|�׵K��C�6;�ƨ��
c��o�u9��;���36^<�Qz`ɱ���qY�J:���(��O�E�&o�u��xu��"��Q������ ���rX���&xbh%�X�ݟ>���%h�:%�z�T������e��z+%ڪ&A�h.!�H�����+��m���# �:�<�3[�zXbZ� ^��E]�ي7�Zf�8�!�� ���t���.)���)������"Uʀ��]��1v�����m6���j�`1���)pv<XWH�"�������RU��!�8bD��{��aL���|�*�h���E�?	S��.��0�B�	V	�����@N� �����u�ˎ�=u�6G��Y��S!h��ay{��c��A�;oی��f�	��C����p�S�ĵU�T$�6G��ݺ������L"_�c6�;х��0pw�ò쥘�t�~�M2����EW3y g=̵xj��lB����zxqx�0���������~�R�V9�z���6�����V�abBW��Na�'�O���G���;5h�b�(��_V�cX��kb�:�z�;���V\-��MGچ��6��oٻ��ս�'p]���p#�.]�*�m����NT��u|,U ��1��f}�9��VG.�,�ߠ�������#q�[gU�O��[��E���1˛��_�'��;J�gs�����/#w�y\�;�ƿ���.a@լ9���Ў��;���N��0�`J��
��>�^�R�����%qn z�;%���{�R\+��I}u�J�F���1Ȗ��?����g��d�P|�&�G�O��q�=��?�y����D�O����+�{��!�<f��A ES=
W'b���p���?~[��-]��{��}C��}k����@��b��*���(l�"�&�4qû1��2UAԃ~�� �3K�_)V5�N$�ţ[����Z��o�*б�3��9P�D[����D ���3Qf����1����RJ1D�ݓ�����!�!'�b����f#M�C8%U�I;�+�j*�9��m.�UtSk�ǣR����'���+�ɒ��~�D��������ꬥ��_��^��4�7�0�����Dw���e��4,/4˲焛O���(i��/��ru`-5c��ri/��N����'�w�(��|�^|�y��oG�ge���YO� �ʐ`��������a}�̚��"�L^����+>�8-/����/@�$.�,�@9�hs���$�8�'�����+8��_�M��u���Y4�>���O�D������puz��l�� �ЍC 7���|�ְ�(��y���æб���T �J�l��p�Z�I�G�����7&Nrm·���֝{�ճ��ә�g*VdA�趡Mؖ9�⥡��+��f����=���ʿU~I�!!k�;��SׄlZW50NM������Z�9�� a�Sb���#�^���ͺ�� �l��Y��	�_�"��5��}�S,�����ų��`3�"�"��̙�Q�L��ԒAD����V7��բ��\hG�/P��(c�)�D���Mٍ�5�U;킩���ˎM�xٕ��Pn.h�;�w�N7+�	�ɰ�F� x] ����P�8��\J�Y��&1��3ܲE@L[	�-����	4�L ��r@{a����J�o콊��D��،|�Y����0�,��1 �7��|ڀ7G�u�q�π��e)%�7��C*�2��P$��;+!��]iQ}[g/>G"2#�ַٌ��N��?p�س����7>�!�+*T�[P�;(�K,':�![�)47�59b��/��%z�P��p�q���` 3�v�w���������WR�K���`\�D���0�X{L���'��6:"�"�
�,��In���ڤ=s��k���E\Y'�$�6m$p�S
���-��vFN�˜�?+��R�&��YͰN�u���������E�����su0kO���ͦ,#�����ow]'>B�X8��%+;OL��)`v���%8e��ٚ3\ �%�C�/�ء��g.�q_g��7���\��A{3���Fd\UM<)6���Vt��@�T3 �nK�zȜ:�2&>T^�@���~�R��>�����l��)�d+��W�5�o�CJ�u�=��.���e�҆��zkѶ���a�l�U�����s��n��b��韢Sn�s��vb#E�UU7��T����4z�(�|b��_Ǐ	�u����I2�xm�T��J)6s�*^����X�'���58lN��T��x�+._Ҭ
��Ѧ(�Nދ�y+�������7&b��z$�0�9uIK��oU�&���y��f;ǡ��������3JsŨ^<����al��i�߃������K�%/;-}����hA^H~��F�a�t�h;�Ì�%AS*_}{�͔񁼳�Dƻ�� PQ@��Ct����+�U���'��F�E3�������%�v�r�)=`g-tّ�ؒh eM�@��F�!ٔ{���jCT�IW��ix��ZY�bs��H�4)Z�@eư&P�Ou��Ҵ�6��<B�@��XGǟR�ul�'��+&��¬�e*;)����5��y�E����i��8����2C��0j�ҦB-�kT�&f�o7��" Ѝ3'~��U���Z��O�A}�c��0}�\(ӳ:�SG�X��~Q�_�,!�f#J�z�9�r��Tl�u�+{��U�q��o�X�0%��ý⁯��
il%��M��j��T
��Y��.Y.�_�,<���ڏ��I��!�Sb�B���9��Mظ#c3�$D���u6H�NnN�^V����.�
����*z�!g_�I2�@1-��v��OW�EF݋�V��(����!���z�G�-��<~	�Z�j6�$��!-Z9� �:IihysgfρPxAY�����]�*�O�0����5��K3!}����D��0ԣN��n���L��;;�����		"�}���9��[9K�ٺĀȵ�>�})Qh<�p�4Es� ��
�/Lo�����eh0�zO BN.�z��OΗm��7)^tۡ��(f�m
�YL�E[J�g�]&�T��'uPv�lnl$!0W�}��bD���~{!0��J4�./�X�XlxV16EB    fa00    2310���;�t�.��r�}\ep�
�)�9Y���']�E+�[6�4f=���M�-�F@u�����J/5Z;2�
��%Z:�#
�4���a�*C��e<�TjW"��e�ig�o�%+2Pn�U^˺�E?�X�J�7�2J�/�$ i���
 �b2q[�gu^G�/a���3�e�`��s��=�=!������a`hI%���x��X���j���؝2)1F�+��5���V�"���K�N9,�o�~L,�h�S<��D��
X�9��g��݊���-'�V����bS-i��	���H��~�JE�2=�ʫ](�Q͕'�s�ӕ�΋� \��)��:7���13?��;�I�GCXL=���]���L��nr�]L�������(��9_DS�4Q�­^�n����U�?�k ��K� ވ�D(��|eFt����ȏ��bR&��h����hrK����w$m���6M:�1�С��)è�p�f�M�m£����2oY����a!�	� 7;s�PG�����4H.�(|�v�撈�Q��f�)��O��� ��6~���k}�t�=��n �p�q4�<_��G�#���l�?�9���8-�q �!t�FG��*��<��/�z���ܵ���V
���U+���܏�^�;{tR�Q�k�ت�w?��R&�w�4!��HgX�8�)�ς:v�3
�ꎫ-Q�����K�ꇚ��3��X<�����*I�
U8y�h�__����f��E���۰s����un|�5:�w�EJ��h��*����&���	�����!}K�|>ɲ������V.����@Y`����q\gA!j�͑?�c��Am��Pz���m�Tԧ��S<y:J=�C�Mq�b`:V|>J�"(}C(KX�Y7�@�K�nB��Sq���$x�$d9X:6�̎��������Fa�sB�x���gJH��1l��\�X��u�	o��G�Օc����W'�G�6V��� n�X�-p�� l'Ѫtr:��|V>�#�N�t�l�#�K�T؉�8*���P�M`�s�GF�KgÎ��!4Ƣ�2_C�w;��\
�8ȹA8;|	,���xh�}��Yc���L��).c�����Օ���R�T�{�ל�q^>:�"ԅ�Զ��h��SG� b���x�׃�&s�n[��-m�[[E\��s�����A]h��Qh��F|�]+�Vy�is�{G��)[U�󜆑"I
�n��(�U�k�ρ@��B���b�e�7e��t���I<�>Q�O���dİJ��!��̘���\��GR���� 7�dJ��M�gN~��i9s�-*sǲ��K0����^�7x+�i�I<�c������"�D$�����4�*�&�j�2���)�yi��k��,K"��p�r��H���M=]��tKW��� n���g^�$���%����[�M�2�y�݆�z�gOܽ��=�My_z{�fH��,`�ӱ[_Չ,��fT���s"e�a�1��SH�����̆���2Zy�I���y�/�N�yr!۽֘X�ɀ�<9K*�/��e'qB��ӭ��T�������]Q�����o���1,��'��ض��Յ���D��yz�*ě�G�͈	}^&_��sX[	�mpMg���N�¢Zpː著ox{�Z������ZK=��~ans�H�*9;���;#삭��^$Cc��i2|���"�:�de�}����������/f�.&4�]���q�,i.x��]b8g��o�Y��vq��nP/G?w��v�m5���x���s�-���E���:״GY��6��^;tK��y-�x�@��!�|ۯ����I�r��H�B����}��ƺ��+�7T��E�̮g,��'�6�ۇoko�;���0$Pz��;���˒�/Df�8�% :��.��n��g���c,�J�U�ɏ/�́/9&AHk��9���֒ ��̺��<z(!���D/f���G��i�XE =6�C��ܣ��ը�G>w�Ѯ"���\K�9��5��k*�`[�d�az���I�@귬$�����@����J�oX��%��>#6;��]��������Ff��lvV�1��(�k�
b板�X��_kD���^J;��*�u���ֺ����PA|zd��5!E�棏L<�S�c�M,��'�gV��6#֫�O8�@��"�ݳ����_�R+6�[����q�h<�mI'�W��T'��{ O�Xw`�).���^�iA �'�N)�O�?���\{��K��*8��Q�?s��61㓒4ԅ��o�T�"Anp%�O�ϛ�IUb��f�c=����5��.VkȔ,�h�}^��o��*2��n��<"+@k~�r$;#��\S	]�HR�Z���w�/{�FH��^��-9E�
�J4��י��+�-��)��^�Ƈlʸ-��?�N��?�46R���S�Z��R֭z��L�K{��/�P��>�YHm[m���1�^���rH�3��FSi*�lA!1��[	P��e��&�m}�?�����Q&��LR{��q��R�hq�57�e�����
��:�eW�N@�Tji°E�������j	r�Z��r��d�om �w{�kW�~�߂J3c��a�hj46�[y���n�o�I�`.Ҍ����9�&��JqE�p홳����xC�EX�*�����8�{ܡ�^����䊱�v�*�-ţ��;!<�3oٟV>�1z�v>9\�[ʏP���S� �7��Ht�I2ϊw*�[,�t�I�s��4������(Sz_/�`�M��@��୧56d{V��YFb	ۯ$FS��o�[W7F�n��O,o���0n�m�&�U�O���A����	�.y��~�W@p�Q���,�(�!�X3��G��6�9B�_����NQ�x�3:Wn��4<*��2t�`&�]��m +��ϑ�r����KO�;���I�F�1���������]Kx��ڽj :.�����?m�����YLKr�N��(J��J���_��XYW6g'/��Gk�+g8����'+������Ӛ�i��Q\a�'�z,"6/F��%���5��y��jƽ��0��b뽉��g������)RV�;��4�M'R���V)A"��K
[	;(E(��W��a��(/ج� ���[$l��q����@��͌O3�*_bL?�`A�A0��E�~����	��)��	�g���!)��^,�})ݤ�[7.��W� ��p��C�{��d�Ӣ����'Ea����̱�,/p�ی�a�}�+YR�"5�iB�g���6'�⛔&�E��n-�O�j���+z���� ���8���r������-_y�^Ϲ�I朠Tc��|�ʾGP�S�`�}w��m���aK�L���9�6�gچ���FT�Ԣ�*�EU#�{鑷��Vل�'sgk�v+o�N0!6x�	ӓT�TA���B�L�����Fq�x����^:��\3�kʘ�ꥩ�1\��ejS��џ{y>�����%L �����CEX0�Msŕn�"����GE?�dN����O�8�1���,x���*��%�?�ܜu���n�X!�}R���\%�"b����$x���	S�v!YB�U�u��X)|������t��u~��׿���γ��iZ�H����壪���-��\�*�
aF�*Ԣ�8��~�9����&.j}��m�[e�*%�שJ�O���l�hRh��8 /��U�������ݧߩȈ�-Y`]s,�n���/���n����*�?����պv5��8&�D_��3wI��D��K�W���+�x��-S�涢��|��e�(��F��$�r���N��z��{����@���=�w.������&��Q2�b�q�lI;�	�(���Y��?�8��jQ�������O*�:�+ $�t��&��I2,%c$Y���\�y]��	Z�c8����ڄ��Y?Z� y�	�A��>�"P�=�Lcd�z��r�����
��H�P�-�R�7�����ƛ�(�o]�5�pU�M�,'�Pp��73�J�����L��4ٙ6���\Ɍ�d3n���c��I~����]$�~���1��3XAB��KPr�˿S�r�2U������� `հn��aʕ���W3����&a����P_-0��c"5��3O�_���!f��O@��m�#-��	�y3�ܩ��M�E'#�P3��u	� Z���C���ă��� ��X�P:�Wa��M���*�>�w���c�"d��v�3$��T��J��a�WD�x'�XL�G��i��*i;���9nm%��F���y�SBN���;�PEUs�!U���<�o�_�֯.���%��31�:��C�e�T�8V��@�~�Fw8@�q)h�j>探iK�$]ZXGP�C@�#��L�^�v���XS�ə��z먕��C��}!>��+f�5DQ�5��'C���L�]����e�L�Djah�}�z��ƌ�?X���b��_�M���?re�`���RqAo�����պT+��|��kXqqM/\�{����Js����M�3��1Nw���&1�sV�6�G}���#�"�jbp����O;�>Eq�m�oM��}�Z�e����,
�-rP�b�<'��~�%_6�m��8�v"�7����K��ݛ|I2�]E�Ou<w�<�r�C����W�����d����6��?r}N��.��8��(8� �q,-N�7��e�u��`�E �;^�z&r�����4۵���oY'6����b�V����M;Lx�]?c %��jeڥM��D���? ���`��n��s0x+���^� �=6y�c�m�
�!��"LWl�S�{���-���Z�����X~^˙�B�*Ԃ�;��m�6`��"*K�4X��RƑ��b���������O-9��Q�|�p@)x�N��򙼢z�I�^/(+��ea�V-�e'M"e�����`���ڌ���]�*��
�6��)/�*��IO����3�M��W�����~�l�s��ݏ�hWu�����w�����V$	���s����Fl��|�ͼ��G��D@�>��8=i;�gǂC�������&����x�ʝ��4��G#����~��-�bh�S�a�����;�>T��49"2Gΐ8X2�#��;�O�H�Ed�;�O�I�'��tɝ>>�9Q�mJ�Ng�[QF�9{3'�k�3�Ok�*=ă�r���m���bMˋ�����H�)���{�m*z&T+*�x>���{!)���]c8M�^�l�8��� l0�Ke�{��5f�]�,eI���`�r���*�$By���� ǯ0�i�ojR'K%���a&��TD�f�lhm>����/ �̮�����}v\J/��.rzPg�I��m	�k���i�k9����'ld��okv,4L�� [#2��b�w3��4��0�xߎVQ*�ܫ]Cu�f�t)X�i���|08��7m����tb��U��y�b]jEU��:u�NG����L˱ռ�<_�С�S\�K��D�HQ��Q��:)�0x]ub�[c#�A ���ʹ�_|!�P���A��*B��K��&Q�TO7Ǎ�%���ψ�4��TUX��5yEc�׋�4��;e�XbH�tU��Q˕Ҟ��8��IK�+�˸����ߠ���{e�����S8@S����X���v��8�9��^���m5�n�`��ؐ��Ba�����7�[�C��0QfL�k���4;��hH娗P\!o�����J\�M�_Hh����E����������K�)��B�8xw�pOEd�M\�l� )eIa/�IM ����^y�j���F��E����kr$p��ϡ���Cۑ
�A%-?�5i6�9���F�.���q�č[ȑ�'��}��R�.t�Q��N������'G����rʹ�g�}->6I긞�X7��
1ԙV1���� ��.���%��	`��}�����T�����ŭ�*��/��K��Mhk���L��{5�8���F�]:�̝Ed���'�,aH�M��յ����ĸ�w��f�T�
�g?���N)kO��F�,._�B[F��n6������U���4ig���>�O��q,3�A7|5fy�6r+�����q��	m�H�]�tۣ�џ�G'�kr�m��%����^��d,��'Y����_)�g2����_��ȫ�3��]GmѠY��hI@Ի��R���f%�S�����$=��)-1(���U4���E[hM���ӧ��F�g�q��H�?�Ɇ����#d��,بDÉ.����DS��֤_��K���yM��s�ˊ�Ot�L���\�s�����+{;8n|�g���ݸ	hI�'���<,I�g���axF }�STn"yDU��XR���7i� h@�N5Ge����;hԯ�y���%��mx4�J���X9e�*���d+|�,v/��i��"�7�8U���G.Q$q�q��51j;�8��i��5~(�3T���<�-�+Z�iէ(�+�9�K�eImf�n�m.�B+wj��R<=}㲄S9vF��NT0�e��j�q;2���@�&��=G�W�`
O6XQ~=)�Mr�[ ������������q��r�����.2N�K���׀�EY����^��I"  ��l�3�Ԃע�4ᎲWB=0x+�0��8�=���5Yg�bk �����]��>�o��HZ� {���������e�Q�i�%���� ��
1ev4�vs�YG��L^n�R�~wl؇�!�F���`�����
)����԰��h�'��lwO�d�(d�=a��#�"sf2&����+�(Y�v9^e�|�J�,�����p�t"��Ԫ(46��ե5byo��4]�2�	�E���z��-�����h�����v�5�Äm@xW��8�_``v�=E��C29��a̅//j>��ze� �Q%.��BZ�c��q�D�]�����@��W�m�#1 	���m}��X��s�M����;qS[e6 �CV���^ U�!D��|/���ȇ~�-q�Xt��Ն�E -&l�y�ߣ�3�]*�����bhr��bW�|�j{�d�g~��"��R�R��ߴ�=�����E������v�:�"�=� ��x�{dOX%��w�_�cJ�t�m����;T�ֶ	桤%���T�øcpуe����yw�����C�갰���t ��L��� 4(����F�����h��ۯ���*d���s�&$=�9j���b�z��J@��6ȈϚ��¦�a��>��B#w]P�RҞ�]�G�lnU&m��=(��	������?t���3R�TX��J�J-|$��;���}�`�����c�����GǍ�j�u~~q������;�oM�<,��IBYim���Ӻ�D��KB nSf� O���*i_�&�$��o����Y���yL]���)țx���|E��5pk�m�;����H|[
57�~8��ؼY,�>�/y�逓{$9أ���b	�v	|��?F���MGv'>c�p��>x���eP�/@Hd��B�����=w��Բ�3���>H4����'�k����T��\C�� ���x�~u�uq�(��$���o��Vո�,��iz����4�G`/`;-Ȼ5��&����(4ו�$�&e������ؙ�#\T֋���֨t<%�~n��e��1���9�&ڊJvL�' �n�����À����z?'�� �i'��#�������'�1YI��Y��F�w�7iH���?ʮ �~�XB�>#������]���,�dabQKj�P5�z�WtEC��sI��X-�n� �AP�譍׎�I���O�D<{h�������k������|p�\��?���5l��J�Y�0�&��/��C ��e=�.�����5�-M5�o>�	j���z1���+�;�o�!�j��+_�&���׷d����$o�E��T���I�3�;v״�R�䈜�.(�K	e�v�H3���$�x����4�����m����Eа�����
�[��!KO?�!&�0^@V1��ȅ�r����&��������Vls�w)Qfd�^����n�Uzv��
\�A�N���z5#^��9��=G��#NL��zT;��<���D�-ҫ9�Y�&&\)tP��~�T��R��X^�\��u��kKT~�'�Ig@3/��$�EÛ�x��_��	����޹r������x���?@����,	��n]۸rS/���9��n�U�?�K���H��"��h4D���2�����]�˅D����~�'aW�jl��*2|�RE�:z��#�}^�t��zY�lY���p��Փ�ݠvƞ���(�����M���9�V褘/���#en����b �-���r ����(iE+��mf�&��>U�IݰP���7��Op���߄!qt�9�wR����Ç@�K�:Fci�11�(1�u�C�K�d���o�8`>����<���$�A����ubb���}wO$�23�Ӂ�]<(�Q�Nx��ZD�81���إ̐sX��EP�	l�>�l�n#��l���lt�j�RR�$��wS�BaG��p���1�"vK]���i�]�v�zҹa��p
)��fZr�cY�	�	�(����1/��E���ꖡ��p7	(bT�*ږ��l�z��e�hk�u�3�(�T��g	�;�nXlxV16EB    fa00    1ee0`eU�)���zO&���������«�\K��8l��V��J�c�U�n=��2����D���c�F�6ws�YW<���6#)�Ib8�+Z����pZ���I��������ܶ��:�xC~�eA	{�][a�`�������'��'Z=C�MT�*'��m=3x9��׈.�����f�.f!�=�Z���P���[�Q���l��>9�Z�m>/�B�ZD�o�<ԥ7j�W�A;n�,h�������gX3h�n<��g�+�����ۂ����tC3�!�zh{��@3%iN��R$�E �d۠���P�f/cNEI.�t䭟����s�e5�����z�Nӧ��{S�� H���ب��z���&�`bN�Mf��z�BL�JC�����S�zK��5�"<-5��_"ٲj���{Y]��o�6�����y�>����s�ũv�G6A�`�xp�K��_�$����&��RJ;�-��B�bz��z�Q�:�h99Q�^l�7^���Һ��D�>t����_���%F���M��-I� | R ����_"�l��F���|�������������P�j���O�����j��zے��v���I4B�Ϊ噪ĘB���αb�T ��:z�(Kk��0�]�)�	��P�>7�Q(8��?`��AYX�A���s񌏧���i/%g�^�9�frl�,�T%��;v�]���7��1d���2ZÎ��w,	�0�v4F����yO!��0SNOsf7p��V�;�>e�)��D���d�1.Z�&T �^U6OaDA������M�@E��9��>�Z��Y�2��D5r����Ƭ	|���&^B�L�C/��	e�J.
 � 0P%���R>e��VW.o?E�<�@Q�U(!�"1�6�� ���6"��:��:'l�<�Pe*[�����
F�0ڴ+>k�fJ>��J��sd��Om	fCRE��u�2��LT�s,�>@Ng2��<,/ֆ�^3G�}Z?�ly��ҍ#n�,P��!��c��z�f/�������j����@��v�^�p`\��Av*ݿ�rz�Y�n�!���3��G�U�<�G:Y~&> V�A��ģ��W�~T�����n1�W�Ҕ��Z�)'��������N@���Ru�3]*HzO��(Ɋ0��	.�4�!�9���P=��"/�]@�_��N9�G살<	�� �ݒ�Iq�-����j5`�>��s��6�nR_�ᦕ�g&�Y�*���v�j���[;�-��/L�};�e��n��!��6�/1����)O-�����_Ċ-�#g \��8��-,�TiMS[���C�QѤ"�Gva�	�:��w.��d%p�ƕ�<�r�u�=U�g�L�l]ɒ���m�������������i���@���� ��%>����Y��/�MN8�@95j>�d���_EO%�~�g:�۬����Y!�*�Rm(�1E�B��3XKz��\�k��XC�}+L���ݣ4�w�T[P6�6�0~�F#خ,�s�����z��h��.��*Q�K�e����ځg��ݱk^-�W� +}Pm��a~Q��Ο�99ߌ��J_�Ak�E�ܖ��N~�[�'	+�SL/��;<O�F�V�ք�ϔ(˾�~Mp1,wʊy�]@��O:�i6b���,���&,=��}r<)+:\j4ɛ]6�;���J+x&nh�8Y�;�.9��@��>�)QB�;�2�l�]���8Dr�g�h�JJ�*7��J�0�f��j�l�@�G�E�Ƚ���E��������t#�Z�%=��q��o��`�Z����oǱ>������a��Q�B�jUd#��W�J�s��U�C�P�P5�.�6�D%x`:h��� ��m�&��9�=�-H����C�=3W�Ҿ^�o���%&f�1���Koh�-~(�p���jPag.���R�6�d:�g�p�Ii+� �3 �,��\s�"��Q� ��i�:�jQ�d�_����P��s�޿C9������J�A��&p����||��}�������)@m�<�0��q�R��Ȣv��PAł:��y#[���D����w�C���?��ւe$��,�G|O9��Ԩ$mV����܂��؝`�r^���J�}1�-����V��_&͞+-ͅ�D���_m����XkgzQ��c�^���<�
`�� �VH�*�R��g�K2�L�_8aI�?og+K��/��p�D1����w�P *����*j���b��5��tdi����*15i.I�rwq������yF%�٣Zڮ��\�6�zu�\���Y�5C�nE�C��hY[XPD�X��Jx;�����,33GC���z�%k����f���)�D5���`_S���
X#�?ޑ(��S���ێ$��&�o]��+1��_Z�A�|��]ro_��Ȓ��ҋ;y� Ȑ�3�$R<N��2�,�X
\�V�[{�б�R4iZ�X}u������=��폺w	��[#���Q�D�Q����z���r^�j�CG�x�/�d���uq܉�E���N�ջ��YX� ��1�x#wT��-���gy$�x��vW�I��+e2�"�Wİ��y���˩}�D�S&�%Q�ނ�T"��/ngi4�r���wݜ���i}4L�&� Rz�~Ǳk�,�(�ٮ9V�u�*;�)	V��h��}�XZWΕx�j։�1������+��E
|⫇�gi~t��L��R���z�I��x^s�]��q|aE�B������~��jB��������MMiY��x�m�2D L�S�f����©{s���̾7�$>1�4��>|< ��$�s�2ۋ<���&  ���x�)�p6Dy��<�_���tT}����e��%e���g�"+��6k�D-����2����<���b�j���ml7#<s�R#������	{'_������mҰ�MQU����6L��,W�Jw,B��Xi� <d5�*~���f���3>^M�mZ����9�%��L2G�զ6�.�����r_8@m�L̓�9��0�JmNW~.jz�xJ�֭&���\6�N���Ж˝]��˻��0��샹f����\y�Y��I�!�+�f�"(��-m?-=;<k�3|��w�|{+x�%�BQ��_�yNH�S��m�z�xй��4���7�F%�0%4��A@�J�E̕��v�z�BȮWf�J7ˠI>�PL��H}[W,	x�O���D���M^���P%��V�h������q�13����55�p�Š�kP�XD�N��������^F�wxF_�v��8_�����d�P���Y7r)��~��j�e�f��7)�Y&����L�U�rs�78��A�L�e�����>u�Gl�z����c@C�K	�d]/��㤵�H����Ռ�ٽ�R��I�(�}OS=��7��?�QO��:cTA@�-�,u��_ht*i:���v2=�6�Ĺe��E��Y��P��2�R%��a�լl���b�5���T6���|`���{�������!�;���,lS�p'��ݼ~e�{~;z|�	�sĖ	�ۋ��я��QR� F�Oq�Q� �	~����:"ay�K#��|��%ф*�"��S����ڽ���-�P%���x�]v*l��7p��궈�a�H���#��q��B3�~!�I��'�X+�zutykj����T�p�E�q�n�� ��p��vr��,َ=�#�AH�čCri	�0�>ٰ�9�I��ӻ˾�������u(Nl~���$���℃f��u!ΡP7�������h�'05��%+96C�
Y1��~���ßy{�F�&��m:��(w~��MQ���Cm��tG�*p��������*99ws�8�YU3�)<��Zu�hH�]qa��#a�~��C*B��4*�V0!,pL����H�h��]e���G���-�Lp�."����0��F�N���)�����#f��:i�uo^Y�l�UAиq��H�{��ym5c8�J@�Ӧi�>�X	��*�cc;A��X�J�̂���>Z��~�X�9/���W'����z����7��;L��6˛�������3dWp��z�d�߃*�Q�-ވ���b�O�D��t���;:��ԮLg]oC\���cu1�A6�8�����(�k���'���O��ȧ ��3��k�*`�Ub�!C��Hd,w}��i�4{����"0\���x�_6���^`��<>ۛ9Μ#R������
U�%;���(��yH��� &>��JΕM*	��n�QKK��_l!�
�|S�������!퍚W����Qr����mU�w�ZNE�x�3����q�5XS�eܣLzEnE���})���� %��'��6<��+c�q�F[�א�:��l?ܞ!��84�hV�I�w�75����`'J����U�5�ªP��?��Skr�q�W9�Q�I�+x �]/��,��w�U����(��b+�Nf�_�D7���C��Ю2x�W����>/�3�i\���O����Q��~�|�<ʨ(f�4J`�:�L�>ɓ�ܐSF�m�����m͠��5�H���Oc�C�_sv�*���q�+�A(=?�^��X�P�LoQh���q���q�&-F)>��Ճ`Q����0��"A�j��/X��h�A�wz����(Q4�I�4���9ր��rh�1B����w��t��UsGY�]���ߡR`�MIW�������'3� ����¬;,l�]G�+�C�]\�;z�C�9���'/�g���#}l'H�T�Z���#��Vr`����u�+~�F`J78駓�d'1�9����w���{�#��׮^G��F��Q$�P_�!�mYH1���\�{���2&�����y
b<�3��[=���t���?�S(��9���/���p���W�����Z�"֩��|bB�gL�gI�n,�I���6S"v�����M1ȶ߽���v���ʮz��v��b��<\��o��n�ƭ��aκo�S�I��)�㤔3]��v���`��s�9.*6�k�,HtK�&�N�ʨ�����Ry��~���.��G�(�s�r��(m�e+�ۡy�62�͐�\(}?��)T��Mf�A|��UP�`L��ZU<=�)U���_K�c�M4�=����s�rb�z�rϑ�DID~���/H}���u������PQ�$ԋ]_�2�r,�7F�b�ܯ��m�u|���w(���7����φ<ʞi?m���V��S�c+tG���]ƛ�x�C�S�c��Ͳ��Tｉ�3le�2�R��jrߋ��Ŷ�0�?�X�R97��a�J� X8;qo���N���u�� |�p�~L>L�`�D��WX]�L��G��GFx�� ;�q�����'��� �@�0�Tt����<)0�U��a����
��ch�S0uj����@�g���$$�E�ih2�zL[��_��^d�V����g���WU"��
���4�/H���8W���Y�~vs��y��G��<>��AOTs�9�� ���_F)3Ͻc��	]L�y��6'�Z9f㒫�OB�:ҁ��g���c� }5|&.cȵ����
�AZN�²��I+K��,��|U��n��'���ԏ��ҋwz���'yH����h�;--���	.A1�ƽ�<�F��"�t�!�I� S�����gB�������a��
���i89�8�s�uXa:o$�?b�����ʐ�5��r����Ѯ�+/A���z�*4��.3S�m�!�=ю	��gB��yp�� �p�kg��|��b�@)��1�����Ii�������W�,>CP��-�����ī�k���N����uz���Ӿ�=H\�����j��r���?�@�.�ˏ�E������J=D9�H�b	>	����9d�FD.j-UKh˗�Dځ|Ɯ�k��
O�����\֘����a~���dM����Z���j;f8*_t��V33�T�F_��W��ax|s��A���q$8TfX�H"�VE�߬ThV&9���Hkߦ 00��d�u�C���̨�S�sT:ވoHd9�됭�0��9�3)!i�W�K��U�$�{�ֱ�5�X9Uv۵���?LD��ׅR͝n��F�a��)�L�w$�ܧ�]9�X��6D����:#��S�mw^����S#�W��&���v���#����>?�N�np ���x��G�E͉~5U�=�_6�9�O��l��ɥ�yP���Y҃E�_VC�s��\�~�@`4a� �įu���c۳���EVנa�g%`K���f~�{Kӱ����h
���p�!9�� �/�#r.#�4�)��z*�(��vsk}�Of��+`����~���FU����oKefY���.)| ���P�VZ���h|"\��:��$$ƣv�+COF�Z��P�
CM:���B\M�5-?�1�����qюK,U�����$b�3rl��\�gv�a�?3[����c��3���@�q����׀g"9�b�y��w�xOT	Ձ�s�xUU����Z67�[V0wr�w}�=�ߦ��Za�Έ/ٶ� ̘($�N�&���`s?�u�mtD�!�$aO��8r-�p���o@k�p�<f�Y�\���
P��j��4�5����t
�\���6�B����e[��j~�U��I"s�d�e�(Z�+���j��'I|��^�5�$*�����Ӿl���S�x������q�fD|'B�Ŋ�	� d�U	
���ɴ>)"J+s�F�6ɰ��B�ڄ�s�W�h� ՉWUD#��#ؾ���J�TM��Ȃ~I�+��s��##I̘�ĳ��5��6
����r=$����K!Kj�k������K�,��"�:�b�Z��;�
hC:sr߾�`��.�r��d։fJAP�a[���W���aw�c�б�p�� ���b"M�5y ������"E;�P��-��f�`�ք�<���g���nk�vph>)hm�$����.k���N'U=����/���4x�������9�>��-��qU��.�Ghq�A��\b�M��T��izz��s��v�)���=���R;з��7w���i<�C�d:�{g�Nƿ%u��*� �����ڸC`fO*�	��G-��"|�>�_���ൃ)�!K|!N+�Y}u*#Ţ�P���N@6p���dt��bJ�i^O�p3k����0�G5�����3�~]�D'�5f�:�V���*tg�Q7������x�)V�[���hR�l2uY��X�U����!d�c�@{�H���ݐj��CQy/���xcw����,^q�E�~]�j]+�K�I85Wd��Q'&�@�ze�T�<h`��t�;�Bt�p���.R7ޖ��I��{5�8,�����p���9���� ����yR̀���L�3�O�oǞj�8��A:�o&�Jl�F��w��g�6��;	��^Rbi���<�lk�����d��:��H��rn�r�P�`�9$S�%�?W"�U���z�k�h�@7,��t����g X�D�譶�[�j���'ִ8b����uE�o��N#WDyWࣞA�_E��9�U�J9��������m�YFdHW�����D*T�)����,��^���� �ˮ�J����|�a�dƽ��p�Œ�S!��X��5=&����vm�g��Oc�t��1�m�"W���������Y	ډ��6.�!�W�O'�ܝ�}���r����n�^���^�p7��x����uf,�E6XlxV16EB    fa00    2250��&4�Ds�On*G�~�������S�xL���Fr�������p0�w�6ݦ�!��S�&z�&9d#]j�Z��@sV�\�[d���펼H���ךD�M,@]W�Y���b����y�J$�-�9��|'�|��Wˈ���d�R�/�P�O9N� ����NV+�g9>Ũ��� ���&pc4&BY	0��K$���;K���b���f�G�������v�˼�,��(m�3z����I�,�y���'��9�'�c:�.�9��V�_f(���6>�oZ���AgZ5���;�}ܺ� +��^�S��m�Z���$��uM&����J&���l0WS~h��&I0&C�]&@�p��*��� $P��6���yK n����AQ�ĤR�컼�Z��Y�h���J��!��M�Eƛ��P�شٷN�W����`�4\񥐚տ;/£n;K�6^c��di/B��͆�I������d���j;P�F���ģ3pcr� �t-)��/q�"���uLջ�2�� ߞ��2�7vXv� ��c2�sV��'���v}��J9aB!UŊ��WŬ��?�f�=6p~�h	)����Z;j[�613`w��':L(��5ʥ��4_]ͼ�4��	d5�-H8)G�r���<�'C沪��*��8p�e�b��FG�,��<yFz_�b۾TF�3R�<:�;'a�j&��R�Ri��G���LY��ܰr�%�iÅ��G�IFԥ&��4z���Â>�� )��<�t�-��.Sۇ���6�U���#�>tt%rd�m�OKBTђ�MĞeWڏ��}?K5~��NMߍr�9h����<6D�q	�z�Ka��M�?�o�j��j�k����g^!���-��`���T�0/��:.0� ���oh5<�:(Մә�:#Q"�r�V�HK���6���=�y��\����i�4xօ��k���˵�o���͖���R+�|���qEИ��6�e��`���/;p,���!}�[�{/D�J�a"����?�X
�K5��G����j�2'��BL{4�1���y~����F[���i��!�kH\mo9����$&PV	�</�miǘ��لP2��*O�b��?�Jrc@�>�LM�SCQq�a�-�����Kx�O��� 瓻�%��՟����؏�U�d��#��߅'�6r�#N ��,Uth�Xa>gt>e��0'Z���E��{�Z[&m��ؖ͏���%�c�_�1m=5$w�R��|���*�]�e.r_�̛�W n-�CSI��WFTJʲJ��:m�ޙ́E�غ�����SC?�ꡯ9��$���aM��Vź�0�����dW�啮^�Kvv ���m%�j�`"1���Ws�>��~ǀw@s�5�JTJ�U�!����E�+֣|]�7�<G�/W�nènJeᤋ4T-^��l���Y�)����qA���*0�o[��)
��k8�Ctѡ�}vۮ���'j�
h�/���ڭ�`���8�VwӼm&���,~��T�Ц��}��iM�l)�Vk��\d��{y�ޞy���Cڹ؏�N6f���5[�\��� !*.�G�۷q%U�͆�$�0���]݃?�n�ܠ���*�n���C�`ۨɵ����0�7��P�@+q{D���%�7��>Rj&�5��,,�S�YBhI@>)�[#�ڹל���,5oWZ�ʆ3eX8<O4������Kڶ�l��يƗb�����7{����-�c����޺E�����#�]x���?�`o���z>�.DFߣ�_QtB�����Oȓ��ӱ��bl��X���]��`�lШ���9.�8*T�|���B5c��������z���^��[w��"J�&��{{��,Q_3��a� z�Y6}���h4D���g�A����](-�^NQ���J\���J�N�dR�����x ����1<�T�	��X'\��SF��1��e��أj�L΍�թM��s���~v5�\�V x~I���W��+ P0��1m��#6�nˆ�/R�0�OV�i�uG�,��ZQ3���}9��`�����ֲ!#�Jr�W!�[^
S���T���C�]��s����/B����@�([���-i�V7=�$A�33~�J���ElD2�&	��'.��Ѐ �Ly/�Z�J�"
��L�gAm���5��'AB��5���+vW᝕�J��2Gy?�j���a�/��s�{�,F��j�4�.z	GT��y�>�;�����X����b��G��\z.Z��d�j���㈏K'v�E4��~�IÕ��0$����P ru��Xȋ�S��:�m1䐟s���@'9
��V!���]��!y�Ju&kJL�vKy��nG�0ⲻ��*�����C��#6�:kic]������o�F[
K���ii��[B�j���J��j�y ޕ�UԀ�j�S�>��d�W�~s5Y~�[gW�I]�_m����.����t%����
�t�ӽ���>�b�[7��[�J�����5� �-,@"� .��5x��5T��&�ם����h�gKl�'�&�:4ҴW��du�G�~X�<�VƮ�^*氻�O����r�l|ؖ��-+�:N�����F��?���5�B��@5��wG�p��Z%K��_G�����Q��`+�
,�8�����DD�BX<�J��	X'��199۵^[�O��b�K��K��0�/�m�]sfi�4�PA��k�[��6&[w�c�rKɗ����(}��Ʃ/���;�T �U ���s�B�RGA��@�fձM����WS� |��w�OJ_�*��j%��ײ��Uդ����٩RC��;�rx�q�H?�E����1�[�(����U�J1�k4�y!�X72����(�;K��*��$������zާwk�©�5[fJ�o��պ��~�M��u;I��d��eBs.��0g���^�+RR*h��Hj7�P���<Y����3���ԪV�	�c��eG�8�������DW�n#�Z7H���;�$c�̃�MGK�4�!���KĔW���Anݪwӈ�c���8"m����}cV������[1V,��P
e#. ���=1�O3D�[�c��y�9Ǒ��ѥ7������oa�>���s�A�b8����+��n���1 ]�`�bB�j�pV�i��	;�Q5R��H�.G�����Oo	C�Bt�q���-!�䵇z;	_D�(q�YG��0��S*?OR��TP���&KD�<@Nh�w�<��=~Ə�3�bJ�z�$YL��΃���;ՁS����,��T������%W�I�|�|X3�D3qI[5L���m�1Hg%,(���h�o��Jy7���2�6����QU��C�C�m��&�?���]!KI�������W�F749��+u�^�Tg\�Ƈ��I��(�l���Hx�`���7`�#c��x�?���f�I����^(N�����Ҩ2�P�){=H�����G Q���a�U���ywJ:Crĵd�ux�?��ХQC��6dّJ��'R�$�d��r@�S(W�E`oY��Lu�_�A�ދ�E��Ր����1�V����8���l_�w'y�7ʆ1��O	�U>��敥�Aj����(�{�H��=�����$6���(�U#E�R�4֪O �#�ZT����W�e��
1��o�S�|�8�H8��%`���w4�(2���hG�+�A,6�l#�V-�@�g��w^	1qS�9���VeJ���+"<A1�SF\\]%��a-9a���7(MZ_.���=/�ĳt��� RK�ZE�R�=Z�*��������LM�vW��Z�" �LuJG0�'�I�����x������R�ryp{�|j7�I����58~m��}���H��`��|IIDYBr$�ȹ��F�����T�#�����R�>/��l}>����>��R��3��1w:��%�B4�m���*7��k����ǀ'扦i������'��	 
?;��7,�ΒEϟ��n�qs�U?�tAq�a7��}�>
����+gbS�	�,�Ƭ�!�GC���}IW��¶�\�o���H^��CL���C����o+�I�+~1}忶b浡|����Cezb�n�Y�ߞ]�:�p�A&���m�4� ���()GL���z���2�+��^y�NWb�%Db�9'���e�g�vq�U�������)ؒ2e� �����?��XPn5��F]��N�}�"^+?�����lz�Vƫ,y�ҷ�>c�u���H�(Mꆙ����6
������>��<?����G@0!�Rp	c�0A��O\5�L_�5lo`��vJX�/�����/]��pU�$� b=�並%$��e�ZE�Ŵ�Px�O-�9R}$�2���ݛe�(�%7��r7㦝R�i|���Ĺ���Xڠ <f�lV4Gp���}v7u:s�j�C�U�u��v�C̬y�j#������Z���HV
��S̫?APݽZc�s��0��~�h7�~]�L�兑�^P=��v��{G���ڍ�:Y����evį�bo.@�Ņ�d��pJ6^�`���g;�Eh��g�ŹT��r��n��X����$!iz��b�4�On>FP�c�P�V¥�Z�C'�'x�E9:l~���"���}��_��Ө�A��'Bf���j��](�GO���{ݝ���5�`�4Ԡn�;NK $)��%�2a���<�k_Is��u'+��cn��˹���ʩ@�T ?�顓�L's��UY������Jt��OC�'�\��>�SF6\�l>���GJ_�߇������/Ԡ��t��x�/:�!'����݊O����<U�s;�v��D��7�#<  R�'��/B���=j5���k�A�O1����lX~�,{5Ţc�	`������&ک�L�
c�We�kM��+����-���L^l�����{��ͻ?m��������� ��g%5Bʛ��W×������@��3V��<f�;C+���W��Ў�fl��XM��VR��d·���Ɋj�Ǘ^��}0VKQ����|���Wǿ�s7��Tɔ��݉�ca�Y�	����42���ok:����H��Z"{��V%�Q���[O66vt�۱�-�<�Ȃ�#��=���_q�(}.����i�:���y�(���a��#rz� p����JV�4���q�U�R��;�A�P �8 �ā���Iw�U?\�1��z
Y~�qV��x�IZj��y�yr!�:Ap7�;��\2�"
�8X^ܠ���/�ٞ#���sz�,1jӆ{����5Ja�L��|�;�8 �E�#63���s.h'Q�D�=}<!<2Ԡ+��:FuC��$����r佛��/5I�0��� <۾��c�*O�iP�����KLP����Т��~���ֹ�&��S�~\s(N��/6�r�K8�m�N�1<���s��z�Uӹ𜗻$[շlM2��)»n��'nP� ������5���LFlv͆ �FlL䔧s�� ����f�u��yO�i���7�JC�5��Y�)����1���n���K欕�Yz�X*3�t$h-1��5L-��Rp���(f9��Td���v�w��^�Ek��^�f燑fY�Su#L�X�[i���^�D~�����xD���`�6�'�ODz��w>>k����vo �������\?�:�O6��Q��[��#�I�Y�Itd���j��	��d��T�X2�*-a����1�Ӈ�ͯ��TT=��Uã57\���n1���j&��������˥с%�L�~�a	L�ΰ��a�t�D ��op�k?'k�B��ؗ� �Qi�i{Bx����ib����}��2��遥���J+"��N����3"*E(���!|ߑ��$��
�'ls:�u~'�j5ks峣���ːl����a�P��g| t� �M�k��q���b�E��Z�{�����J��.�i��q]n�t$C��l4��d�a�jԍ���U���rm��v����yg��jH��#���"(��5�Ӗ|A���vVd�x�KC�f����Fp�#F;jBRv���-:zn�{�3��e@�� �`��S�Eb=��U1��۶ѱR�Y��:Cآx���&y禤�AMxlG�6WCW�)��
��׼��JAğLo}�(��������j4��ӈ&S�yj��n����t�	e�:�M�M�L����p��|�a��b��𹑽[u�@�Jw�\v���:�논���9A���
��2�_!n
T�c�`��fa��	�v���J����M�)�vm�}�λi�V���n3{!�\�m��m\�� ��PkVT籪�<�OmZ�N[ی�4N�e�كa��qj`��8��9g������6�Hòx��}�E<�3V��#�~k:ʠ�D=�@g�vǦ��i���c����%�^Ҏr�Ę�A4c���pS)6���)�V*��;���mϴ����6��s-��")Ɩ?049��z�נ`󈗴mw<�{ԯ5��˧��!�qsM&N�i����2J�yڌg�pf���sl�m]Ge��	��Yh9��|�!��`uVr�X�z<e�"2_�S���==z����ߌT�:��Py�[��˱�^ #�<��<o(���s	g��扶�x<���3 *TC���H��>)cu�0y���7qQ��_�1�p|nSU���Yݢ�	�V(2�pt�0�N?wr���j��!W��v�4zq�e��7�(/)[�9��=��F� nWd9 Bc �#�#�J�,t�P��1FvQ��_ ���'=�f�Iպ�}DL=��R�$G�9/8?�:+_d&@��$���3'(0-M�X��Ԥup<.X��T��9�D?�!}z:?��8Ta(v��~|CH��f�,s�qi�!�h�����-�0Y%)��������85�&z�2��,��'��@jû���Kn��'˲bEܠ~��x��lX���;�	'��gO�@���%�_��q���SE(��gy*m�+N>%2}������`�!���cw�Ɛ=&��f�0|�g�.]�`�\�sJ�m�t>&	k��'݂|��>��y��lpl��1�S������K���28ic!'�N@P���z�K���y�TQ~�֨W��}�O�\ۿ�<���Z�~Ǡ������.��t�H�p���n,e�E�g�7Q�5X��zG"?��]Lj&NbT*
?����a7���L����|�5P��?m���Q�Ǆ��d�P�6�Շ_va���� �C���A/6�p3�"�p����d�hU�K��ͱ���͗�+%3n�ar����F��d3�9ຏ����V�=Y)���d�H /�_s�g����+�w�A�0F�ؾ�Z��G)�e�I��u/��z{���fP	ާ��QY5��-��6W����&���;��*�V������s��P$�kGF�P���`{��g;�U�:��x���߉ >�]D[ �����Nn^��(��;��Y����8�2f���{!�����6c�9ԷlI�}��q�&H��,΁JxU<D���>:Ln�YVxghgЫa�Y�����W�G�fxR�Ĳ��x�lF?���Q�ڮ�[��?�D
�A��!|k����P�%5j�����Ƿ�M߈k��D
��$)�l���Z׎,��~�R���R�{�ȅ�״ i.�%��'G�~�h��~=��5���$o�:�m��$����f(Y�#2���ib�+�,n�Ȅ;a�{�^k{h�w&�zը�,�=O�<,���m�����V)��y�zƵ���Nؒ���e�����w��.���.��*ë?�M�Yهn���1���;X���� >���)ݎ�˜c�F���W ��/_gU$���ߨA-����1��]��¨0z���U;�[�ER�0x:�h\^m�HR�[�/��
��x��2Ldhg($.o葁��~���
�H��I�wʢ�����2|���H�&�烤��A���WPh��>��e)Yb.��aO~6�#D�ɚ�F��Yt��C����Co���WE��f�%���&�/*�Oߝ\�V��[��m s�%/��̢|�q^):eL�!����V[�v$��`�= ��c� �����,������{^�
�G
��,_��}�r��`c��k�Sڄ�;������������e�5��6s�>�,eS���g-ss2; ��&H[� �" <����[�i�prV���v�u#������cj�|J)Az����wײ���s #Ұ9�_�#j�ϱ#���b`��ŋTW�+|r>l��I��&�G�Q���U��=T�Z��8f�7Lۏ��kZG'�%������(�d��\j*+��RwiG�	*O���h𦗧0\ �$	>pK��Z��B,I�ٳ%�ʜ�kk�����x�Y�'e�i��o��&{٠Nx�n�]�R>��U�E9����z�����H���� ��>�H�,]Q�y���
&��y���w#�j�%8��d7m���>�K_�
 �!٢g�c9yg�n�tn��f�Y��~vL�4����gi(M�p�����t��\z5�3�Kd���q����F��ްay���
ד}�Ƞ�%5A�i��jײ���Χ���XlxV16EB    fa00    14e0®SGL�&��`/��KHr� ����zϧ��}�eS�Ś����{I���)�R0/�����^YLWqZ���f}0��M���e�ke-��Q|�}ѥ���m�uw�����.�'�c����?���
�}<�Ph�����ǋk�a��!YP�����P�Q4�埁��R̜��eR�����,b�J/�&���K��V���1)nq�����Ģ���n��c�P�8L��g"�9�)�8$��UGNF�f�]���a��=A�ɯ�r�����J�����N�=��'OB��ۘ!��E��Z��@�fj.�52̌2�w�mOٹ�p�͹��Rߞ���t��L�}�xN�:���VdS0cڢ/�F{35�QN4��0]Y�#��bt�慭�D��d&-�4fJ��CJ����.�ۚ��1a	���U7�<ԥ{9\��	q�2��:�bI�{��q�ߞ
��ӺQ7+p��o
�4*t�"Y	��rm*����$��sg��Q�~�_@e~d/��6�Z�f��?Lgw��8QӼ�ꪎ-����H����|��q�e����fj0��hEb�|����S�B�l_��<o�O�-�������d�JV�ӹy~͊M���M]��Ho��xү3��APGVv,hy� Tu0�t[?���-0�G>����J��	,x��t���z����R�M�)�ޑҸ���٦ ����[��z�5��[j)Bv��hF�-£����7�'�7�F\=��F4��%K����|��ɀ�(:i�:�:Ø�^���R�L'{��&��c ӟ9S��H80l�k�K��t���<j��|�Rpqu!%�t_�Y�#���B�r�=�v%{��$BX�|f]s�tn�]�M- ����9�q�\��-o��P�����eJ\YL@�0ŶT�����x�]gMN����#��ᕼ�>�u�ں���4��A�&�����|B����止�"���t1v�͋�㓐5���Ê�'Y������t����0��eF:q+�&��~�! ���NO�;�)���G��;G
�7S���H��$W�������+�r4�ܽ[�{��.�'Fm��YYe�f�PH �h���ɲ�5������ag���d5�ˉ�.DG������:ǿt���oŀf��a������~���~ϲ�f�b�v!Å(��=ұ��pW�&�/7ħ+��l�~x��
ߑ��:��.��L��xF,�������`�u����/]v�%߰�|/<T��jw`�>�a�o���B�j9kno����[����F���R� ���^o�{�
���K��$�W_��Ԓ���߾m=N�����xR!���N�?�& 7��.���:8�����U�~'��Z,����)�c�:7��ŉ�O�؇?��\Ou�X&��������^�^��W���M�Wh_J�Z�$u����H���Y��������z�}E�*{���gJkj��]T[�1P����:d��S*�@� 7�3����1G
�{��D�' �;�n��i���r��oiI��j�F��VB�fZ�}�P'Kq�˷M��� ��a^-�
OZ+��T�o����=���qq�j�9B:�>F�u={����������Ŷ�+���j��$A���D��?� ��Ԑ���i��Vz�h\�w�ԫ&���ښ{Ew �`;tu$��T�`lGy�@��˻�(��#�a�-}�8ws-H�.�.Xˎ���g��܄M�y��j���4+�eɊ �݌&�p���G�(�%�\>�,�S��2�a$�Z:V4��F
�����g���
�dֵ���g�X��İ�e9Wp���><���<7�����OC �u��������8��RQ�yh�~��$.2�Gp�����p)�m`������Ĳ�2m��h�����P�t]}b66{�o�A���@·(o]��,����3�B2��Pr��p.��������~��$��>$�R��]��7�#�pl��H�rh���6�o=��9�{J7z���G�	(��%}1�SpI�t� �s��r�@3[���^As|������gw��4�G����L��B��mj�����Q�z�h(���i�p�P�]�܏����ꐓ}��;��P�ŗ��~s�NP�	�~l�������7H��Qc���A�DvB��2�ׂao~�l�S��U���,��j��ʆ���{JǞ�|���璓�mP_P@���zx�����NE�ķ�:�"��TD�(�\�J�_B�q��+��I���z<Buf,���Q�փ�RR�X|��.�c���T�c�����sw�"襩�{��a73�c�t� �"��gΤ*�R�Gnt2S�/�h��X�	��-�4�c	W�s����2�E<�;#���f�sh\S��Ш[�	,t?������4�N�źAX{�󂙒!��b���}VkeW��1L��!�.����6HJ��ߎs �]�$����>'��~,�3A��y���:�&~���^���(�?�S@�O[yrY�77w�دۗ���-gH�.45A�;b�K��ecqv�J2��P!݉m_pR�����RSeӳ��.�v�VbL�,�v/�{*܈�<�.9�J���v&����~�;�X|[=�?�k��|���1�$�T�SK栎%_\%;[�<S2D��{�g@���Ƭx�v�X�%�Ii�&���c�+s$R�5�`�O��� (R貚�մQ>c/Q� �$w��=��K�DF禍��溡9�*�V��nJ�0l:�U�d@���
� O$p�����DQ�y�_t.9���n��4���W�����Y͏2�i� i��GEf�^�SP�� R#�o%�QC����ĸ`�q�Iw�^6"~���ǘ��3~�3�~�$�\��3��p����v�b Tu�!>a񼖫�=�M���!�y�~5M-̗��2�?᭢�)�%�\Qб�}���#��gN}����1�����X�
Y-��"�M�X�O��qi�Ʃ;`9l�{��ې�z���w.
߸}1�ZGK���ݬ�����bXZ:EU�ɾP#?���0T �DE�
��{?i6��&�MQ�!/�a@6�D�O�>z�1<;u�dGT���-�\s�P��5����r�k0���r/V�e"�E�ʻ��~�}�g�:@��¼m1S�CS+'�BjP?�>�$�J�ExLLR�t�¶G_*((Zƒ
]�/1�._��ޛ��n��������j����f6�LFFۆa %a��K�����]�8��!��]
d{�9%�]��n�E�"���-&�	��z���^��g�����C0��d�O"�d���c;],�⣘���������9���,53Hu>�ć�ȯ��	%��,��	�+8�aL��c{�:�B�����(6|g�ђ5�`���O�i-	�,^�4��X��qSE�HM��P�P��Z��5Xr�����7IUR��i��%I�{|�~��a̧��)���q�� qw��Tu�`�K�A`Hi��f�K]B�韙���E���G��u�p�U�C{�����p�H݇������[����8�q�k�֣��|C�$҉��g�a�� ݊T�F�٫l�ėz���ﳩff���Q�[A�Xn� ��\�����CF���D�Sl�3�R� ψ��d�$^���U��Τ��-�m��R�tX���F��&�&��4&�؍\����+W
���dG-\Y�^+*�"�R�.�	|��]����^V4?�"w����r�γ܀�la��t�%F$J2ď��"�T���%�r<�� �D��C������kb�Y�g�',�޶'1�!�\$���o�c����	��?�b��������*j�P�����:O}�sKli�4�AP�>0��"){���B�/��)�X~�3s��	� o��6%���u�y�Wշ�d��'p�h��!�q����P-C���׿�I�ۃ�)�ߺ8)�RS��D��/��N�9ƵD[����t�c�R��4������T����+�V�H�=H��"_A��FŘ��b��J���No�q;l�"��ٳD��qy-*u�"0��R�P5�*�}F�������g���pn�/F�b۷���D��7j�;�樚��u"Dk�����Sj@��K��s8�����E��c��CvӾϕ��c)6#h1��Ț^�pą)�Y��T~"�/s�*^�{{��[Q�$:C�e�H������r���󷇺1�lFg�������<�O��N&)�b�{v�m��'��Q9���r#�Wٖ�k� ��/#9Z������~h�"��.���f%�o���_�P�Cj���L>,&��1l�V�e�!�P6�K�}����U"|���;�	�|���4KP�;���7L4|Ϋ�;�������q���;��V�9y̾IJ6��][x}�ʮ{W��X�U���ⴡ��!X��g���ξ�c��x~n� �iѻ�Z[� ��
������~E�&;�����d�uZ?�<��|������<��D�����zg�ʆ�Y*�ī2��3J�i_d�/Q�s�~�)��FI��i���#n�5]����$�T�ؙ/e�W��z{�2��x���Zo
��IP9�J��� ���c�B�`��-���ޔ"V\��=���Y��:���5���P����$`w9�q�C.xs���I'�CG��~|���t��~�	�Sι���=�+�K�Y��MȟDX�D�Ł�i�7�歉3�G�	�R�|'F:oV7j����~+�[���DT H��=��φ�A_�m�� ���茁�BM��Q�E�N|B3fj�y���N7u<����3��|��G���i���]1��=C�/�1Do;��P'���r���Q�Gg{�~�`��}�x(��P�+�3@A!�Y�����N�y�{�sL��)�f���ŭwBX�_�p���dB�=	9����݉������o.!���q�8]������T�'�J��r�WKU�1%�v�i�Ba�;y$� k��I-����~�� WHl��&�9X6�c����6�JK��!/o]Ӏ?���v�zw�?��U-y@vo��`�C?j�E�nO�Vg`�7�?%N��̞ɀ���E0��!b�n��E�V��<G��&_���5�P�/lҥǯ�ss`
a���l;�@ˈ�'B)M�!#~���V5�Y0b���i��h�XlxV16EB    fa00     e40�`5H��=pW)\�~%�)xQ&��0�TH�\�>�n�g�u�?.k@:p��I�LI� �<����7�/�	��LS�~{p� ���vՈ�{
�����+k#�PL�l�\��q��D�{ ;D�bE�e~�O��YG�*����w��)A��"�vc�\�7���y򸷶�_ɴT^�J��UL<�P̖R@�RX`	���G�R;�K?oL:29s;�h}�����w�7���KZX��q��
��5��K"��1�i)H;*��e�@a���?���*��}�������$���?f$%���EZ��97�6bi�@������H�q��rw�W{��De^_\YT�ֲ��t��ՠ:
\�!Z,��:j���=�4y�~�A8ҿ�F�S�OY5�6����f��'q"��6���3M�;FZ)�p�/�GB�6\&�T�y?	ۼ���{f�i�xIZ�Nv�5<Y��p�&8O�����_(�H'���7�Md�ҜP�c���0�X��n�
J��4��HL4�\�8޽2�?������OT�eW5}24a~a��9w_Vc�má�Ĕ��[�Z�oX�O�kY���JX�����!�Y�2��/�=JE��	��%�`�	i��8[-�!�R�	n�`gqe��m�VU����t�R轀4�6����w��@��Q5�	X�����f�9D ��&�9�Uƕ���{�u)����la�C���~��Ww4���qgE��W���گ7��ڎ��k]_Հ��r��=aDe�0�u�J�����,^�&A��fav�x�"��,�.V��Y�+\��6nN��R�vj�S�<S_]���r��ܿ�J)�ex�E�~2��	�z�b�9j�C��~_Mz��}߂-�.l�`��V,�=�ڗ�[��'^�i�>�aDd'�Xi��I+r�;����G��S�Z������W���He�+�_Et1����+�N<�^�~�q��?o%N�ڨj)񗊇K��xb�vS!��3z�#5�/�3S��{x[��I5�YN�� ����9�A���َwO���@4Q�� J���v�)5f�[F��Y�y���Z��HǷ��VJ4{��A�L���3�F�_������J1��J��Y���[�
=ՌԴ����N���.���HH�ﴫaD��� җ���p����,���2�wv|���i����[_Lv�=�Yz!P�4����H�H5K���|��U�����5�8l�t�v��L���D�;�|Uj��mPբ�i^T�_������LD-u4�ToL������ל0����k����c)�|�g8ʑ�� k>E�U�f(V�DR���Iv|�kVԡ��Vi+�Ť��O9�����<�_E1��7�%�EZ&n��@:}�&��1L��9*�Po�x��7	��z<v��o�e����h^�%Em��ňT�l��e���]��<�P}�ߝ�<�Zy�<RE�V�&�:�D�R<�g��h�E�f7��55���C���	>\�ш�dV��Q�^�^'��#�Ä��5��@Kõ�@�G�/��*�uCɬ/N���J�\p�Q
�T�����òm�.��h�q�	G�����~��'���&��ipHU��Î���"�N�>9�b�ޭ[M�A�M� ����0^�f�G��+4䖱͊��P�5~#E��ё,�=��b4~`�I���&6�N�<�N�\�[�����a������^�Vv���ӏ���t����uMs�ʭ�"��	�-��0x�ώD׍���h�ut8�}��/��kkr�b����i|�7�wB=2�m�bof��kx۟"
(�(ڗ��z��U���]|�D��+���Vԝ'�F���L4�??� �]q���C,u��h��&ϳU�5m�@.b�l�_������.��GW�B�@�N��ꮻ��\3���.uDF|���K07N�"CyQ����V��~zJD��Q9�����=i��u��D�@ׅW�R� ,4"���X�`��r� $�S��t�~G���9J�	���	���^���(Da�� 
��3z�����[Q��E)�Jj��d((}��v�}���R<o�z�#��sC���~1,Af�咅 ���k�/����!��\�*}a�E�.Y�Xd�'���Bi!@�.��<���a��
DY.�!w�^.VӻP{ˠa�]Oy}ӊ�
q��,�1C*q?|A�Y�ؕ��&��Y� �����v`
o�����Z�}����+�(�P���_�ձ5����l��0��A�B|� ��	Eg$�*1�d�V"�cu@�L?��̷
�����_���6�������W�N�k>>���w�]��-��vӋ͆�b���m�c$��ۊ�I*�O�ޱ��I]0�x2��FM�ӂ����k!~�z�Η����☩��=�B�@�tjM���[���r�;2�~"N�f&W�X�B��g���N[ao��N糞J��Ae?/�����}Y�(]i����F,�� ��r~4Ȫ*�"xi=q4�4�;�$�@8-ə����o�k�����#2*LF/�Cj7{�E�]~$DK�W�~j1b�1p�2	���hsY��S�]|#���nz�s'���u�s�w���R�h!�T����+�ˌږ��p$����`il�`��s?Ê��D#H#y&b\K높�k>�JC�;d�&�)ݯ��LH�����a���+�҇d(��!\T���.{�f|�&5`�XC�	�����,.wmrF����BO�37G��j���eu*G��%�QQ�M�g�S��H3e1y�Pe=�#��>?ә�0��*Â��U��D����ѐb�+F��G��,��I�g1\m/��W�sSO����>��b �~��຺Gŭ�5HOw��S���yS"$��۟;���N� ��~��u+��ee����r�$�"�	5��V��ǵ����̉���W����q (�$|��r嶢t��S�=����,F�h+R�����ie{d^m�v�(�N�2/I�n�+1lH����=��i1�uXY��������
�M����Y����?cə�g�0!O�
L٫
;�����琊�&�I�b�uU���ۚ�1#�����Dy>�}1�G1<��}�+�@��$j��� �e�L&�_�t����[�/�C6�YzB�ڎV�jt���,'Ύɥg�c]-m��Ԭ�m�9@: @�Т�ݰz|?(��c����?�T�r�����<��%�C��?х<(�B�ı�K7T���nL��Ό.ۜ�mD��y�h�pA>`޷%:�%��_�`�_H���ob5�J�#;�f�n�FӨ[�����KBAڨ����w�k'��Z~c۟��ߗ�(���� ڔ�N�8n����Q��vJ���i���B!��J��y��ËY�+M�Q�R����|�-̣�iz�2W8��%]E?1y�N>φ���?�y��H	j|-<��1 a>�kҗ?̝⢽�����:C���c��`o	-x��t�ȼ\{E|�X�.j�\����:t�o������1U?"���&��s��Z+���zA����Ss��#�Jbى8P�s��/��Ӎ+�K�XlxV16EB    fa00     ff0�%O��(.p f��Rt�$�p�F=��k&[�(V��!"U��G-��L蛕H��a]�?�)�x�.K-���z�c]��iA���i�>�����RysV�]���ҸJ8L�|p�m�D��0b�>�7Ȏ����T$f���Z��NI^G�ŷ�>�� 9�}V�h�8^2��GZ���h>�>�^�|i��^ǵ_�6��#��NEIⴹ���I�% VA��D�� �Yp��C�{��e�}���Δ��x��A m+U׹Dؿ9��O%�I�Pg����)о�������(�Ĉ��G�|;bs����qP>��%z�A�&��y����C��2`gh�˫���42k`��8���A�g8w�����M��B/�q؀�����!K����J�l�7b96#��H��ƙ�!�]wy9{�-:\��K.���TY�m�VRL�����ߥ�F�!]����~+7�v���,i�(l/���?+?s����.�W��3����o��(8�X���>�����>8�����e%Ջ��@q�5���������ҝT�ߜVmi%���B�ua��'{��D�����&̢D"��Ek��C�N��uQ�?����Is���C>XxV������^�7�������r���2��Oq�Qa��HC���ƌ�1����i��� �.G�C�<Vq��d�V��
����ܧ�Z��i=숇d�W�
�`�i;�8A�%���5��L x��zzǃ��y��<I5N�"�����"����A��������/Zc�wz��]\9�(#����F?���x��à�+�S����t��dV!��t�#�t/�0��F ޸F�nʛ�����0�0u������r�mdH$(n�`���x'��Fn�+vH�l~F����Rl4�k��[\�hq��uh�U��êG��@v�>�>��}+�4���::����䓜S���هt�� B����|"mjQ�|_��W�u*�Пȹ�W0?��@�(M����01�W�۬������s��X�S k!⚂3�k����������]��jޑo�<AQ5�󻠪�%Mt7�ag.��#�'W��y�xt+�Y����&�G��Ѝ b���2�:UQ;I��@�@��'əKIny�ͼP��c���**�U��
b"��_+�,�q��J���)�nb:O~ΡKd��A�������#"W��CM�VK��8�+�9��#ձ!��;C�oV�	�-d�ǈ��R���l�Q�5�6�� Úb?Կu�O�f��Y���0��ߔ��	�cn1	�'�Nc�|��uO;�������6SЯ�QJ���XvoK����j��^%A�>I�p�2*��{5V1b�2r�E��8/� ���&LO"����L��Qu-�9��Ĝ�x�~Z,�Z�;Ӳ��X*��4��
z���(M��4�ͅ:4�X���$R�����j�l� ��Hl�1�h����S<\؈��ou,����1�uY��%�v�X]����;�������K�?-�F%;���rq�bBff!��UL��,EDN����=6�8���%�D�=^G�#k`�C/�͚�F�'�
)�lcH��	t�t�<x��q�;>�$���g�PY�a��B=���W�;en+��]���L)/�(/�_�)�ϥ/+�����OC��Ӳ����-�G/��i��v2e2K�lQ��|'��ϛ� `k|ish�7�W*�Y+�
��Q�����Lū�䟔����1����'I�{�j*��h���@���l��V�w{ݭ{�[�&����{��<oCQ��F"j4���Kơ	];u��R@�o�`�m�ߺ�q���o)0B�� u��y#Y�$����h��T�o�V}4��i����p��U�\^J>��p�/�|ί���̥��4P7�_E ���x�(̻g��r�;6j��F�9�f���}��=i��'��Z>�g�����~���l�:��FfZ~���4�4��?�D���oQ��ٴ1i_1_�0�*�,����m+mNU|�a��f^�f}`�Y��}�n�8�!p#�����b�֛Z%�I����5���9O����UC\p��r��V	�!��o|�/۹��im5Ќ�t7`��y�`]�8CWOHEd��Sx+Uh��3�H�c������2��qaQ���䖜v88���/���ŕ�}W�e{���&Uf��5>�j���W�Y�B@Q!D5��Fa#v��7ҳ��D���0� ���[ݤ���넲�'���S�i~����=WVڲ�vG`�x:V2�θ�1۔ל�ȧ���\�� �c�w5���qc �@����mހm��}o*%+�uc�\���ڵ-HG�A�l����ݛ�V���kc�R
e�XJ��g��͎�3Jj��[�xDǷ�Lő�@��l$,V4��h��8Z�e��N�8���o!�Ky�ì��yi���xL�V| SFP�WU�ˠJ����+��)"�M�,�ԍ�+�Z��Ri��O�����DI�>�3�� ��
Acw@�d��	l~m����'.d��P�ńF�*mP�vA��(v��9Xd�!���Xs�]}�0��@ܢ�Xq������������Y!�b�c�-Z5y� ��-L��=x��v�6�2*�n���WF�;V8�wY��ܫ���異��2MB�{.�X�=�YI�k��U����:JM;���/B�Z�Y�h��V�@J�����i�ˢK�]���r��m�}d�"�]'�Da����ܾ P��78WN�t�2�n��M���bpj\z�Wc(�^����-��3F"|�qA 9�Ǡ7���}�$<ig!�k���X��K_�稣�/r)]6���z��9o�zJ�����1�:E9MR�1�H1��L�;U���y���T�I�DG1V�z�Yt��`�{J#����/���%ͩ\�_9ā�2O�pt
p���� ���GJ�>hė�����t�?����^�7���񽫻Y��Ii�����E_�KU�T�JNQ ��a?��gA�mbx��W��%�s/S0�� s&\����cK�t`��^d��6asA���E&�U���X��{��_��H?+�	�!��`S���Q<"��v#W�^%�}&0Ⱥn�m^�ۤ�"k�-�R���L-�E��'^T1#\�5����d�=���e����r���L�ǭ6\�h����TH0��+8j��;�.��Y��C�9EgO/f��Ahe�u�~?�� �y� ���^��r�b:=���y����׀�t������j�"�T]=	�z�,�����Z�eK��]H6���\�>j=]OT@:��.�l��d�$�b�a�[�}��ّ*Vv0L��
�HE�W^=+��Xmx�̽��|N�#q�������Bls�����~k��v�qz^�__	��"��̀���;'n�|¨}��C�Y#��{]����{]��p9q-�e �x7��֖�3�.�J9C*.BH����Ǐ�+;�X��;H4}��5�,.��Z��|?�m&����wh����K<��s��%\1��B��O0�+���~Qď�Df|�?�J�qR@^����"����K��P�~��ͣ���ѹ�?�p�W�p�6_���蓗8������r}�J�֬G��S�'j[=�M�6V����_��}�h�*�-�}���*�i�ƈL��{ԥ:�.e�[0��.�{���n��R�SV��#���z(ͩ�\��v!�FdՑũ�ݱ']�)���ȵL����-�:��QBŽ�:3a��3y�����X��ʟ��������Tܘ�߼���|czC�Y�ɶ��MA2�/������C$W��}�fM�����K oA�B�ڮVN��X�_
aN��n_`���sY���+��|��8&����t���ȯH�Z���{��"{@4ࡐV�Ǳ�.�j�s��inM�`����B	'/d�k��A�	�u�'�m8׻GX"8��^���W���@��BAXlxV16EB    fa00     b20ft�H��x;;EJ��lJvɨ���d!i$ș�vگ�ψ	��r��aZH?��/C���%����0�ڕtc��]'0���0t����A��ٱ� ��0�[@ۏU �Q���BV�*1��ے:����Z�-<Q5�/����Z����&��}`uv9"Qj�:�8��_���kl�p���tN�n���kW��PDmioe�W^z|����a7Ƅ�|V/�)H�g�*f?UUϱ���t$�
� 7��1�hN4�a�����Q�+�T��HJ��Y����`��r���e��N�{;�Y`,���>'�?UI��o���|Ax�����0���ձwU�g���5V�	�zNϦ(���ˆ����c?��`�����֟���C�$-�W��We�//��e�CX7�$~��qr�
�&��
����ݓ]jF'�jKa�&��i'�ݳ�0]�yRT��CK�c�[�T�f�E���#R�n����7�:���l6��#(k�,�;UAkmcB�}�� b��Řz�&��wѣ6/[�5�s�~��f>GyYG/��ɿ�r �uV�\�����'6�`�
� �|'T�aW��?8�E��i��⢰���Z�{Р;���J����@��W 7k���j'J���Bl����e��F ��� ��8i�]u�����f�OQ�Ԛ��jC�eN0���0�7Z��Q ���	�Ȼ.�Ѽ9��
�O�'��|'�I��x7�[����s ��@DH�Bq35��v�ڶ��aZ�t�,u�@+���!��=��g~"�Dы���f�O�%���V�M�x�X�(C������5��+V���)"�Z"-D�[c�����KaP��,����U�m��a�O�P��诊���4"�4�JZ��Vs��dg/<չܛZ��_�xaäƾ�}Q�z&��te)#�\؄��ٰ��ŗ��$�t�K�~[��x��p�!:��V�>�t�� �!/y�t�f���ϫkT5�|�c��2�u>|�AOBܳ�,�t��N�68M��$̄)�s/\Db���%������S7S�X�M�B�2����n�����
oz���+m��Uc�N�^�.�e��WY�׵�cWT�M���TNu�#O��"�+��Ns������6�V��WL:�-�'z$*ⱴ�h�'�+�LUN�y�������'t'�����q�GuK���_`�Z��>��_}�)�|��7]N��߿�����WÈ��"zK|��, r��Y8hc��9�^��$�ߎd���j�l�#p�Ƶ	7Ѣ��^Ū�IԴ�f�jA��J����K��ΗJԶ��!��	?���2p�ιT�g�W�zGnV��;,}�������ڲ�c3�ݲ۰�;�����u�mE��[AU��R��g����T�޵Ud��&"�[���ߞ��u����[Q��+ax����oW�c���G��\���c9
�v{G9�QO��
|qY�"We +�����E�I?�Iz�w��̛n'�Z��B�1��"Km�z�u��V�ڣo��o��U_F��!��!���s}+#J>SPu'��(��͉���׽ d�}hq�O����^}���7�����²���1x��˂'dY�k���9�E`v�x�r?Z�8���c����\�ZSz.	ŧ6�q��l!�Suu��b� ����=
�Q��:�F�0�1?ETH�tۥ�8٩���>H�ȱ0Y38�����Z�p�N��}�PO���R�C��i��G�?����-�,�A"֒��|O�F�9dz#!:E{Rk6*;?m~�jP��1y�,�^ZpV���(	��m�|g �Nv�u�d��k���^2J�Bͱ��a_�(��r��iL�W
������8��CHi=���.��ІĿ���2r(�;�E��7�L��>J�Ҙ����%�#�	�����i�Ϭ�>��S^� �v�guķ���:2M�4h;g�Sr�a�m֛��������z�#;�I�R���`��i�m�����1�8�?��ߑw��'O@��OV����bjaS��7,��A�Mv�;q`3z����<"{�|�M׊1�k
V���CA~ z*��Wk�_��5B��W�����'�L$>�4>7Q}^ӒE�m�k9Ve���C*�R9g�XbxΗR���	�e��O!MV;X;ksk�}��'W&�x�0����8�R~�`��ۗ�Frs�73y��Ky۠t#D�[���/UI婱��� �<@�r�����|g�NR���WN�I���*M�4x�4�	�W7Kb�J3q��0�:z]�*cV4�?s(�L��R�4�
J
�i�8��S�������)x�Yi�v#��T���v�ׇ#��9�Al�M}3�^�JA٧m���l�4�s��ѯ0�I� ���$�0�>P�C�ع�B�uQ��Ng3u=AG��Ngi��moUG�=�j�HQ{�(E��i�K0;<jx�G@~&&0�2G��͆Y�Tk;�P�w3>*=��ż&!�L�0 �)�Ba��Xb�~AlovJs���Y�i]C�`�~�rW�(���n�=�#�A/ɓy���i�Sn�&�bu���᧪�$O��-�&�K�Rt�;_ɷ��?#i�E;s��ϗ��Mqs����˰,��X䋴c�ݹ���1��\NX0a��he�2�S��u�F�K�Ey��U%mQE�-�Ċ=x=p��͑�[�$3��'VB����;���q+\b{��j��<G|r�`z��%�.=+7y�����j@���,R[�ELX&��8�&���ڪKO�ȁם���g$H�rpXlxV16EB    fa00    19a0����\6�+6�g&m��Y��˵a���@M��o������s����(�)5�(����'L7��u�jJUUNi�&����X�p�3Dz16t�Vt���(4wo=��,y��Ѫ6q�1(+��z?�k1t[��_�I
	f����*��_�.����
�'�j����a���[�fc�lss
T�0��P �w�l�����5b�q-��X�"�>��go�⨻4�����"�l� @sDގR/�CEp4~�R
L�
h��W���.C�#�$a�_��|�~ڪoh��.�i�e�zM�?��u��#��N����JH&���5����릘�:�cJ-!�Kp�~�b�8ƕx�$��m������d#NKp�M
���:�1tD�9�VL��ͮ��2��.R���.<�s�(�
V�AD_�?�Ԁ���V��L���rK:ۙ��Ap���$��7:�#\BB����(#�#��(��^�ْ�]-��j��xq�k�O@���1����(���)I���C���&��+�<F"�to,*'Jб�<��'�,g$���ב�ƪ�)���d×�cb�����|9A�K�`w���;3�J�_b�ȉ�Y�-ho'�;=�.�Az��(U{W&&;���-��AKj��PE�d���E��U&J~]wA��4A���޽����Y|�	����)�B�uq_ڳ����)�6��,��깥���N���Pd����S���*I�I��-&��@,�!MBG�B��S9�x-�h�3�ky��W�sa�TR�ܽ����pwo ����E�j�8�<��v�<!�f��_ޘ�S�n����Y0 ��u���`?��tx}�tމ�zI�,B��X�`�EFHb�E�B'����	y���8>E�	h�)����I)hܢ���3�@�u����J�c��&���V���Gy�� �VL	�l��F*M������)�4�6}J�߃�����Cc��nr�5�b-e�<sccPѷ�ҟ���$���3���Ь%J��_te�0���Äya��j��7��Z�@=0x��kH�m1�.�a�*�e����?��a��1��;��O��j~��E����.3�5�`e�([��pzx[����!��ߏ��rW�24��X�3ፉA~�f{���|��w���g9x�%��>	����<��W��1�/�䩅��������p=<�H�t�h���/Md�C�N��F�-�E��Fqǟ/�'�x߆��lF$EC�&����ÿ���r	�}f��8�]s���@cQ9"��Ld�<�^ӱٷ��O�e��-��
�ʐ��u��ne�c�A��7��g��K�ѷ�i�"�?^s�Ds�����g\S��vD�¤ݼe�Ć�w�{���JS������5�Ab�7UL�)I>j`�������Y�LX�`�����N���"�Y����ձsp3�kbe�r��>��^nǒ���mK\+��R����|� z/������J���jK�:�z%�%F�Ť�f1$�^x����)�d�r�<��m�J�%V�ДiE��@�a�hA�y�|��0ȕ;T�O��+gQ�-P�c��Nh��"=Lҳl"/U	����U�ѕ  "�����3޻b;-�) '���$?H��p,�4��F|�d�
͊��|�q�~��\�1�;�$��E
���q42h�jMt���1�~lr�����U�_إC���x�:{$=�x���`�5�����ߜU{# U�^]a�`�J&=���eؠI�K����T�FJ&tXa�IҡHl��M���颻mX讍k�q
�[B�CFr�^��X�~ �y�*U�UA��A���oˣE�T�v6��9\`ow�x��ٸ�NH�:A������b������T��}�ܷ�N/�2�J$��oZ&1�f�wCB��u3�@�S&Y��!<���g�8�����ab��m"g�"�f<S�ԙ^ʥ��n�5��A���v"����B��fo��G>@a�qQ��:��I�:0��J�~���m;O0O��R�ֺji�É��Ik����o�<�%��#�T>8�tV�u�I�0��h�
K� ���dH�(��5���%L�H��H�y!��4����F��e3�-@%�&������n`ʏG�2���K��êH��%�igQ#��^�qp�(=�p�h� �%�iԓ�-���Tz�a�ˋ*/��H�=��Q|rK�y�T���~C�06��Vb��W��:��  ���x��j�J����0́Yay�/l
E>��Ʌ5��v�"����_XX���#p����M�gV���2��R� �3ub{%`���މhZDM�4�(h�#���y��(��-ۥ���������!�8�x��/L�Ff�r���"]H�^��"=�N�̔��>Y0��[�A�&�Js��K�#2xn�U����w����+'��WC��`!����G�\mg�tĆ�P������0�Y83��Oz�z�k�2����x��j?E�?���]���2�u���A�nB0����y�\ķ ���9�2!Nؒ�S�3\��hR�G��g�s� =�>�����LjN'G1*�\���<��9����:#:�I��J(
$�ַ��UE~�Ad�����Qx&�A�5���H(HM��Q=5>�5�\��� P�Јau<��E�p{���C/�*��dLGB4�s�=J��b�Jԡ��=q�j�����3(���t��FU�����ŅnLAN�*��Mm�IZ���v���[����i U.�=�U���I� �7��z*Ѿ��X����gX���8p��]B��Q[��
�f�U�UHS}:S���6�s����Y�60�T�q�S�����5=��F��%lN��<�$i
^�"a	�c3��
+��d��t��|��׃��H�cb�����&ҿ|>G����~����1.�>�*C����
H��P�k��%�,#�ŕ�$��?���y_w�ޖ�J��9DŽ�m 6�)�6�M�{���=8�/��9`�X:*Z���CsF/wp+���ڷ�*L�~���x��GEy�E���IfZ�~;ʬ9*�����!��,���<�i�7!���n/�/o d`K������VC�iR��v���6*����C�~���ط�5t"�FIv�ң�M� _�*�#A&�j	b��K �_ifO�ř��*�=�����h�"e2}Hڠ2����$�e4�S����yF�7;�]����03���@��+T�����p.�٪`�jqBY�>���~m���;��Kb<��*��
�l�y�[
��-`�ƙ�C�A�j;1ׄ�s�e�#�f�%���i�\�N�ti�g:�z�5���O��m��C'�_���(pn7�:H^"~WM�@�=���V.	��h��V=c����BnjR����Vޱ�\ZR\s�$Y��V�~�YR��*���$;GgRgB2��܌�x�5�(�]
�Mmo�C�W��=|�WL$���b���>e��&�0��!���$�4zw2�i�u3��r������/����:ͭ��j��?��T�a$jK��{����"H��ꆾ�}�����O���7�q���q��U�;`�$��c=���B��o��]�bw�&t�u���c�����쏎���f�BA�-�*"?�p�F�x����Abj���:@s��T�mߊAP�|w�з�nl~Ca0��%c��LmmZ���ɉx�5YF���sU	�2������X�ѓ�������_���|��]vo=�yA�h���<_�('oTW��u\K��r/�O�E�R�skʩ����3�3��3�o	1��b��Konh�VC��:_�u���l�ߢ8p`�-M^�#5ɾ���1�+.����\����w"
����#�*Uk!��5t{��м��ޫ�����!�� �ǈ*+Y&J�#�ss.[[�5l9����;�1<i�pr^���%�Y�(�� �[
<1��5��2�n��D+�����%�B�9���������n��V�9�1��=e��/��=���9� ��\���-P�cu��ϊ�-�	�1P0�-�~��i����!,]��P�3����9s(�ny d�=�؇r��@��Wo�r~{�;`ÒA���������\ s��s��QY:8�������?x�ִ����'*�)��a:-t9��,xA��.��}�ʺ(G�9��T��86��R�AչMq�uvX�q	�SqQ�V������5ip�$��Y �q�(�v�f�H)�N�ݔs�w}�t�`�m���J��\��ks���B�)'m��^�ˊЎ/L�}"QEΕ�w�K?�F�v�����:���:aAI���z}��b�u�-��>���^R����,��m#D�:��*�l�Ԃ5rG��l��P-su΍[$�7ke�.��-�:pn[G���D�Ȧ�l���� +x�>����O%:��۬pI�dP�G;�֞X.ov{)nt���'Ǫ�=��a�����c�Ѻ�J�Z #mȢ�	?�l0�U ������PN�{`7�X��} ,��>���.G0	_�UIu|ihf��5�dJ��D���(�̛S�}8)(��w)p�J%�`�I*�I�g�L�P@
<�GEỒO��c����BU�v���b��0b�7iH;��P1}�D�I�I��ϪIЉl� uNV
����E^��EW�	!2��n=۵����a��ͬT����*C�b(=�i��>+�S_ ��Fp��fv��B�w�ԛ�En����p�7�Y셞��Eܟy�#Tv��e�@��w/Jx �+]i+�!�$c�U�ڪ{��y�u���s>�v��º�U�k�r&+ιM��x�����S����J���I;��c؇x�Շ
m7G��Ȩ�zj�����|�m���=br+o��r��O��"W�d���R<?hKh�D bL�SiR��PUp���F�u�Y�~6hP��\���?�y��}�8~�(�̳)�!��M��x�P�,��bۙ1G@����;�­e�I��,-��xF:U��'?����K��}���i&���|Pˣ��g��+[pF\�{���P
*s�W����%y���zp[��jC5���u��:��5���ݥ����@�8e��1�Fy������}8q�����5����Z�ʖ G�c�sy��Y�1��ݫJ1������~y��,�z σW �k��'�"6azLL����q��V8���F�&/a�G4݆�͔��U�f?I��ɖmp�R�4��*�f"R�2vk�I�lb6`_#�h���c�JrdI�\\Ƽ����s�����)�x��p�Y�bV~>zQ|��j������G��Wi�#pɾ�ؘ�|"���|��!���N ���_ �gS�7�c���_/ۅ�уr�l���,O��Ɯ0����-������`8b�a��Jb�<�WX+��H�P��~���O
�ܧ��h[w�(���r	�uw�(%<k�pǼ9��@�j;�|�?��w79[
�]�#�-@����aڶ�7|��w/}#�xǺK��7�UO���}3��q��o"����{I����Rc�T�;#�;vR�i��k�#j��=J'Fc�����/<F������a>���,іy�yǘK�k��/sy�.^�]0~#풉�-�/��%�&��G��-��:�?<�*~�h68��Mo��� e���z����dGL�9*����
��QC����\mn����ß�&�sw=��wf��3=�9%�r���C�yf�Rc��oPӎ� ��oz��*�����ɧ�c4����}�[�O��')0 �/@�t�E\�]�����2��[~�Ş�����4�%Kՠ墳�V��R+�Ŕ��q���6�%�W���
��.U�!�Ce�e9�SxS�� �A��+sp���(�I� `0��Z�E�p��l�O-m���M��+��З�H&���;$���f��aq~�1U�0�)fn�
r�|��B�}ȍm-����E�&�xB��Lu��*�����Gn&\�g>����@Y��A���8S�?f�!�/�2�	�%��
y"xf�FH�&~��Z���N&)�%���l����qJ)ͧBSH���2���mE[�}I4���N7��GX��mJ{����@C��ryu����Ti�t�8�{��#������E?�k��<9U��2�yK�J7g�lD`��} 0���
�Ͽ�*���3�?f�mӀ�gʇ}a���FJ���d�u#���(J������p�L�>Zh(��� @6����H����أ���#Re�s[�,i�Jr����Y�f����qQL�X@ ���1e���ޜ��(K#���lg	������_1��[��b�_ŻՎ�XlxV16EB    fa00    1f50��ޑU���ݶ[�}8�v�G�\�*=q��G[��}N�m��6����-�W��:r��ڍ��Q�}+A�l��q��+k�х�+�>Υ�	7��:���̱���gz0�j<�Hk=��㋔-?���A@W�ƙeH��FԾ*����wZ��&7�a{Ķ�K��+�W@w�Us�c��_�^�j��ba)P�{�Z#9��!nxm�!H�a�8Ee�1�#� #�G����ڿ� ���H
@ڵ��ِ��̋��_����gg���e"��hu����uA ����cԒ�Mb���Tb `JiJ�]��	�u�� G�Y&>�����p�$ɵ�j�ӌ�>�X�9xi�
df� X�I�߄+���+���͝I��}�bZ�x�O��P[v�y�|�Y�fw+Qc�L/([���Ō�,Mц6��yN{;ZR �`Rmm�T���Q.�Oں̄I��5��c�Sw�@mq�@KM��N���H��K�b]a�F�ڢ�
x�W�N$��_��3-ғ�]��ɐ�:��3�9Z���R4hՈZ�#�<e_�_��K:6k�1��7��K��?l�Y�na���V�����h�k���(TW�L:�7��n����p��Q(�Pԣ�V�'�v���)��|ւ �&{�Y�Z˱w�BO�
sB�熙w�������g�qn:d� 4*r�(��A`?���>e���U��K�i��, !ֲ;7��k�YX�K�N��K��?5���lHv1��_�a�Q=�%��A����V���FM8Uc��D�7V�͇����m�`t�1�w
r@W�m0T�������ݬ�G���UF�
|�D}�x����8U�ϻK����i�6�e�Y�}Yj�OE��JĪ�cٖld�a`��f&ZR�kSI�c�����s�ɾ"��²�癑_��N3��ka�B0�����V�T4�2���[��:�i��d����w,8v֑�u��AI�3G.3�9�>+�e�=Q#��3M�L]a��������1��|m�k�>�IcUl)N��0�va��:<&���:�o�����Ky8�%��>B���)��*������$�����F��7H̽%.�LZ�k��b�@���2�Rq�ɕ�-W�ΰG�o�Q�C9 v���z��^^{�V2"�c�_�*�Is3��#�����P��׋�5����Cv�/�>�X�} +�.NI��燜�����e�y���X1���恑�;�3+�
��E"�%}K������NN�ЃZ��,�i����*c����f�|�Y���˿�[)�X�pb<�J8��.�?�g��ಎN$N<�|��U�T�5�[��쬫��0���+�(��AT�89�ꭥ-�n�w.D���`_G��"���b^��6Ou��p�����»��B�'m~9	z��)��&��h_Y����@�R�ӞHw��`_$bHʒxC>4MWm|�Q}���F��Er4�]�G;۟1W:�Yȧ�^7��_�Rp�Q
���kt�
1vy9�@RN��8�a5o�s�+�����;9��|ze�DڄrJ+�b��o��;C��P�5�oP�\���bK���������!e'F�9-�^^��ED��y����3��З<niİ�1���������y�~;Ư�IOB��P�#_�� <��~����t��g=���l�qܖUd�C�ܑ�Zn�H)��'ru�ر ?����eA�Lv2�e����`��m�����B��.?[K��l�X~F�r�$���T��-ő�&��� �۔@��N�@��s�'��dn "G$M0�P1c�1�}�#�#���k>R��������#:��G��	���Z	1*Vgp�m�W��_��&���(
�3�L/�2df|��� WQ���I�!�'Eb��)t�꩚���ޥIRbE��g�|?^2�"VJe'�~2� K7T�u��uԂ��-�E�	��4�a��#�\����'LھU�B3x�#Oܷܷ�#�s��ZU�h�$
򚶻�s&S*�����܀ K5��C���w����H�F"�� ?ISTR}��}�;�6�+Z�e�Kj�٤'�Y�����J�QXO�S��$�t��Q�a�J-��qp�����J΃?�6���w�~OyT�Eq9��(�:ްoǊ�S�ye,�c�743m,�kB7�ij���i>	��+O�H�7�
VP	@P��8V�>6�k��V�0:�s$�l�qb�R���� 5\���J�l�+�� ׅ M
ǧT1������d>M���h|
����O���4&��25����]��y�}'����-[�;�T�d�T$�v��8�9���ܰsbm�2h'%J"����3GۑN�*B���Z��=�+�PZ{<�54@�,����b���8�%3#R��R��oBst��1s��J@�u %�f�wP�����8M��oĕ3�1��0U���J�,�~��˽!� ��3ږ�����ʓ�j�y����Ȫ,��9��q�C�����ߌnd=` �qIH��.}D鱌	�����;\@U������h�=�&؁_��P��X$:u~���1!?pT�4e^��95hr�H��V1���g�.�<��T]����$�;F^I$��-ݛ ��!�r%��ҊP��t��a��DNwg��/eGg�R�}�&�}��<�K���R����Jh̻���ȺgXT�I��o5������G4ϻ�y��4>�Ǵ�37��S!�d�>���`M��20p�dE�F�8��?��9�����᠓oQb�/|�L�|��@��f���� �32C��aL�B�&<�s&�b c��<�yQ/��0����ᡒ5��d���7 �;�[:�!��4���޶�s]|�F��P�5,q�&A�5	"Z����c�N�����82���_X��-���ç�9	����L\��~�z�[�����wZ)i����J�~��Jp�[�RT]N�=Z�!���ng�˺]�DxRe������u'@j���ߘ-����Ye�H��J綻�Ů���Ν��S�.�6��>�Ov�+D�JH����vf5�=���r*V>��F
	CǕ���$U�g6�e�гQ���>�}d���U~���߬U��gs���sZ�;K���:3��  �'��}	�'\/�,4�-4t�����M"��W��qe�C$wo��t�����~�j��u�[�r�X��f��'0[
7X�o�).��rcL&���1�q�sxnv�,���pDJ���݈����^?�Kǋ�ޣ���ϢLJɲ������Q �_W�ě�
#l-!�B#�N�Q+F�x &{��@��~=)����v>�8���FH�ɉC0�>[2�[>���t���;؉ަ\�x��=~� �q{�weD6_��d4!��~�$,aj��^� ��d\f��p�1h��E���:�^��}Nt��z���6�X)"D��Ծ��l�Б�Y~a`%�X՝�af�Va4�f��auצr$��y4��#c����"#�2	�y�#�ڍ��0�]gO���� �sT�8>��U�]&@��� `P���J�߬��O==�� 3�����������<B����6�����y��^$cq��)с������{�́x�ߥu��i�}"��LVW��z+��� �C�;1�f]������;@r��;AO@�kЋ��r�8�Y C�z�8��#�(����f�e�,;#ٗ��
B����w�o��i�Yo~v�r�?�6r��ѩ�Ѕ���L, ͟�����Jz�
a޲6z��hn��{R���m<��pe�;��V��L
�+&<	"�����xV��P�5ھ�{m�R ޣ�İ�c��c�8 �	g�l�~�&����3��$���\����)y����(>�qL#�vƉ1��2V?K	c��}��� FW�I�U]�%�����̕Y&.�\���SI��"IZ����q��ߒ_����p���z�D�3Sq"���h�(3�ߟg��~���Ǣ�����<dl�Kp7��u>�6zrR����a|��LJ3������Y����'�����]�%�N(��I+��^a(&���t���w����J[�qL������x�mRg>���XF�h>�v@�~�����m��V���9���f�ʉ�0��Cͪ��i%&ڒ}Ԍ��ZjF�"�|d��͖ b)?��%��y"`��q�
d�L�j�\����"�)�#G���2o+��D8���ͻ�@��q�?��ܲ��3r⊂�rC����)���$Yk�Df�Xd���RH�n0P����`N�>�ۿŋ���Ob�|&n} �HTġh{i:�����;��為�g��ӗn��R�-IR8���2�8���{���"H����;� ������Gt�z�4���� ��)T���������n?"-c�����ﵥ�Jf1��!c�&���"��'������8+@���D@i@}����=,�w]�QhX�(]h����1���n��+��2��� }X'���T�9�x�y�
W1������#m���f���R��=Љ�0���q4��k�<���a�8�:�,������Ye�*�*f�����^:�@���6&P�����_�ł�/�Q�x���S�h�6�ލe�s7I�p�:�c���	�~��t��H���X]��j��xt?:�kp�]��(��g87u���K����6I�����V���M�f3�����u��Y���T��GE �X���)���������˖�{689�A�;i��{bΨ��Le$�f�H����A�\5��;͊�a��3����3[W�*���DB�t�����~R6���FQ<_����qP��TB��H"�k�E�^@/y���9��p�%PY;Y"���g��e�J�7ȼ�bm~�9�c%��J.��3/t�;���F"�|�1�)����e �!�H5��4,�����G$�@�aĶ#�tJԑ�!�6��}�Le^�vrQ�Qg�gr1;0L�0[^�Zɕ�x���</bӯB�ܛ�����W�;��yÐ(ua�8�H�Z��v�Q�������d�0��W��qd}�i���f�Oqrd/���S�=,#4�X�0���q�6T��!�]��"Zs�d��@��$&--�;5����G�ڶ�:��]�؞s�XD�Ns�l�95FY98c���1O�O��*t����cD��{�#�f�ſ �R��v.9�b����u�i.��.���Ȳ���ٮ�[+n$iY�36��b���S�>"Dm�!��e�9@�� c���gs��"+"\�䪅 i�E`�Z�B)�3w�a��� �Ό9v`c��?�T����@!LU��{gt'+{3����$�5i�"o�㱽0���B؄�="�|�KL�m�p��đ�����h�u�K�Q�|3�2�4�'�X��e/����|��%��! �8K�de�8�9iX�X�0٨D��j���w��
(ff�*���+k�c�t�j.4��8/�=��Au8|�`���qWs����Iu���Pd0���ū�OM�~��+/��bV��:����M]H�%���a2Tc���_$�)�4J^�6����[�B���b�l�c�BR���oꎿ49�`b5̿}=�IGz�	��3�8�C7ZK�� ��f]$'&8u��Y��jꙪ{'Q_����S��TD!}��)�v�e��]�� Wþ�K��p�e�{��y���g�W�{�6�W�ܳ�yg���G�(�D�?$���+At��З4+:��̓�-\=��j�6@})K=�$�ܕr������+Kb'�| �"�!��[m�0������"}�܇��H.w~��p��S��4+h��[�ڵ��Rx0	�1����i��<���jo��9
���dy��A{�vf�y��[�
v
Xl�+;+๤B%�QY)#mŮR[�p�����.�@^`��J��3����/٧�p[Ⱥ�;Jqw鯝1�B�dђ~�R��%nQB�Ţ�a7��\�.�B�+R�]UVۚ���b!�-����~Oacz�x�vʱw(Oƿ�<+
C�"�c�r�y�08Pl���3)��Y�r�����3«�D�>3	Qm�&EαǬ4?��~�r!	��F+]�Q�3����_9���Z���.�v	�;iL��=ɯ��@�U�2�y�>�vv)P��@���S�	�dNU|���y��֑�y�gi�59b�i��&��sǱÍ�\�ʈ>bcM�V5��΀���%����2m�*�(/c��a�!���`�9-�A^�<]��v}�T�B����O�(EP�<��S
T���#:����s(n��OW�V����H�3v�� �P�MO�C������[|?�5��y'
P(��3�m�s�˖�Ɨ|�>M�H��,��w���n�J]7A9P<nv����2��|���)�����TS�QP
\W�:puu�稰�m5��ph����$��;g��ȁ�_����V
F���gu��z����=�ןƅ-M�'|��w'�;�{��L�d*CM��C��&_���Բ�O��v�[>t8��OZ?�U�Y���.�\t^�m�_xb�"K�k��y���g������q��)��G��J#0�56�g"|�����Y�N^��`�WT=2_= h���!Оs"/H|$x)��h����{�*�g?�а�My��S-��ώT�My�j�m"RƮ� ��m,�t�0����o)��
��2�Z�u�)�ƅt`�}
Χ����'�-�W�ݾ�m�'�I���i��(�0�f��0�{��w��A�"5|���#F��O����A�>2��2�e���̂o9ŗ6m[�2�S
-� 2eG�G�I��ʝM,������_>�ՔZ_�'~4�i)���gs�.?$$�$�#�M��.H��S@Pc�nG� ������+����$+:)k�6D�6'K���ڌ�A	@�gc+���+�姾@\��Q10�zx`F��d�-1Cx�@v����ŞY�ɝ$L��0>���_Y%;{�{!���-L:
)���.�j��
�ٛ'J�����OC��c�~pv}m���[:�b�M\>��S�e��m�Z�n4��"ٓՔ3i�qw�*��cv�^T*ݱ�,Nۇ��d�<}�0�4�R��Z�e�rje�Q	� �w��/]��&�$Z^�I+�2ץ��D����k	��QCmT�\�+hЂ&��Ӌ��c�·�G_Wc�ϋ���5�J��<��J�G9P�G��!���us?㫥s� ;m��wA|ެ4%����MZ	Y(�Cm����c���LYdd0֊+�ABR��#�1i�h/-�=�{�h����o��r��$�"��jIrz�� �m���L.���@��i�����%i}A��D~]�kO�A�HSCމa1��­��ׄ�k�sL�h�3�ÊR�7qEZy�4��0�Q�	������
�����.����W����A�l�t�>�
��ǟ�Qh�[}ORK���uB==��f=���f��9���:.��s����e2����e��>_~�G	����|J�p��_
ʠ3�=�2;�k�@17��hh�˓Xk�OL��7~Վ��J1���;�zˊM��XG O%�e~��-�es�qzv�j앝����&AZr�t|�7���ś����S�.���V;} ��^t�x��vp��������F�u�&�˦E`��ǁ�v�WD!Ǌ z[yi�ln�r��\u��X����R2%�;m'�E��]VN ��s-�zJ��',�lj��J�#B����3�(ɔ-�@�$gsV�NA�"l�g�{4�b[��<�C�ɴN2d�_�v`$-��h�i$L]%L?�S9�w:q��A�7	;إ|�
	oh?Hm�}gFHl�q�W��XlxV16EB    fa00    1890���$w^z���� iE��uh ��=�ȉ��|�.J���Y��uHܐd�v3FOH�����&l��XB��]����"����D�_�Mh!��^�Zjw�PF�� �!���&��c�������Q3B4���|�@��T(N��D��;����������l��i�&�f�������$�7����^�RhM'�&w2���3��Z��L�̻��^�GĲYlQ�ə����Y� ����Y>|?Kq�c��E"��]���=FH>�������Ve#)2�g��Zx���7Trn]�������i{f���)�C�*�A��*�{����k���a�	�a$���-����+����ϔ�ޗ�f�ݛn z�y4X��kR%NDX�	�>]�+LJe�*F��r\�]�(*��[����ߍRYK���z��>!��v�P���H��m��÷�����o1�χ���
}l-�o��G��ʩ��;��S�lL�4��,�U�樯�z��#l����:l�R�0�iw�y҂��]z�D���	_�n�# �x���es|*�R����p���W����Ȋf&���D�`��槦h��(]�W��po�Y���$���ކ��ˁ�T�z{��$�3��������%�)'�1	��]&m��řx�+Ӛb��1�^�Wj��F�y?�n�@,%��5�ޓRHM,��4��g�?5�X���[��򌝠�~����}��t���bD��� �l�t�R�:A�ũ�A[�N@�����K+{@�9ۓ�|�� �x�[ۦv>b]�ٜ������^�����x�X4Y�6=۷X,����#�e+�(m�26�x2ChCbeA����:'m���Tdi�s ��H0%�؀���IꘅV�Nh�וlg�JA��شs;
� �����̊T�B�/��]s� Y���H��oh��pd*mp$1�Ȉ&4�b$
*u��a���8龪��!�J�Uj�xdEi|�^%��;�~<�����h���l�DR:h0[0��#�|�.t�h�r�����6w4?P����/�?�0s���-b�� 5���xg����? �Ϻ����f��5�{v)������ՊN�~�q�����H������a�R)h3���V��Z+����Llbޜ\o|8���͵aֽ�c��A
HEc�%
�ܵ��N�t4��n��l�(�N��2�>���]����s-��) F���O���,�k���B�[7����2�*�� 4lq���ٮ���������g���ְp�+!1\���ȥ�w��G�{|���+e����u��h��f��[�=�����g��,m\��^h�^Ox�!��o:1-��#��5����|xG)OeI�XW��-�q7���&mO�Fx%��^��'{���!  81D�a�0�$C~K�8@��T���($4U��P�a���R�j�d�Α]/�J���@�x�k��Nv��lfOGyGy32���et�N)�s�tv�1�[!0+V&��ܮ�fwkyK�.���,�wi��hBb�fp/�pcP�t��P�A��D�����=/t�}P�d����:�0b�q;�o/�u�t�u8�?������-�@��k&��� ��l��<+Q �y��[V���#�9�-��H�n�k��@H�Z �U�i����A ���mI������	9(��}�-�?Z(���{��W�'b�fW�Ud.9����,��U@J�t�F����l�J�)m�؅��Jb>WT3$˶?��I��;���.���2��С�
��%��/7��R�Sb��#�|��oy����.�ן�[0N�I���w��{�iY
�JF9�Y2b,�<����(�q�a�C_=�������֛'�����A˘^�^�}/�է�1�j�t�0�oYd���<i7O�ۀ�,��B5�`Ok��E�֔�B>c���P<Hp�C�j�����6I�4�� #�Ze��H=��i�o�,2�O&�eSqǻ�O"`q�`�����ki��%�k��c��i�#0.	YѪ��;M���ۭm1�ևr�'�a%|�N}������%�ƈ�n ua��鈽�3Sύfܲ�C��䩲������ڷoG���_���<��<����`����P�����˼ا7�D�� �؜�z���Y9a�H�y>a�Ø�AF���頼�GS��� ��>m0�hMw+��s9߅�Ȳ��M.�)����+^��S>�U`�"� �Q�/�����b��N��T�[� �8�"#�E2��W\XD
f+E��^��NBNs�E�T�R�70�m�E2J��s��������>�i
Fw���9��e1^��|/�j^.6Kj���r�d[�|$�1��U5�T�9�,D�tZ�� �p=Ew�~`R�S��OqW���!Q�ZYDM��5�)=7ٸr�kw�8(:��ৌc�p�%orL�M��QX3�#�i�P�5�j�S�vL�zN�d�d2���L�����-A� ��ƽ� �\�85�ӄ�GT�뗔݊A&N��D��s�[�߾��bvy{��	#GHF�]T�܋��.|�$�V������`h�6_��+�:��;�K59�����ؒ\e`�?3��8_d�s��p��	������*�1-Wg\"�?��М�N |�9�{����N^�swIfM��~F5�`��8�&��0Z^T��]d��!8�g��{M ��/�A����{Y��7;3ILh"f��-�&����f����ʅ�(l�>���5$��2�Һ��I��Ð"i���J�4k��w��~��t>G���D����*�x�y�����VǾpx,Ge��T��F����AK�A�=��ki�E]�Q�r�}C(%���Ɂ��2a�H�o���� &<���:
�t�^F�|1�ϬkST�2Ҏ�����1~�,�:���������Rnt�U��&����_���_D�~�\#��ю���%�y�;�镼"C�]�g2��$.�ApF��Sco�9[Q�5�Q�z����v�$�QT�xi�5��'`yffm�x���I���Y��5�:�?�V�D�i�8��xO�qһ�fvk�a��F���FxGu���q�)#λb�ou��p�`;�	~/Y43��!� n�o��>�Fu!��c���B͎D�Nd3����K��9w*����)�������K� $ � ?9��\,ry���qu4���Ӿ8[U��[���8�hK�zt1+�IeJGs�����C�B��'\rEⵕ�ՆW��p �ss����G�WK
<]�3��{�ǭ�s@�p΀+��ӽ6vd�iQ߿��+fO���Ȉ/�����i �k2s�jB���������\�^��|�nk[��\�����F�U*{
wR�՞`�����v�~oI��n�NI
� m�ӝ&���� i�!>�u�GP�V��VmN�Z`�6ni��t���8�8�7[�t�Q�{��t�Oቑ�7����2pH��L�^@"AX�/^��y�tdls�
���?L.�$�dv
|�[	��0|�%���b�	<���I>�4"���Qɮoз�By�W4%XTU�(���	X4�˓ Ꝣ�����-��/��ǆ*�2}�7������.7x�>e�!+ZJt�P�I��c���$Z�E�@-S��E�^��8[�%���0�/�@�z��2��e��!����7t
�Z�+j96�
�F[
�I:DN1Mj[f������dB���u��G��[Z);����Z(N��$|�/_������|�:I�^Ј=����Q��`^ˋ�/"�c#>���(��e�&���V�!Y��f�E�b4$4x�`�y̴
����y(�]�!L���{?�ˈM��!��]����C�F�7$�aO�@	�f�^�=��H%Y-0倨�ˤ��ox��|dӠ��G�f��[�o��rnS�4�2;��7}��uRy�Q�k�G 'v�٘G,�oU�t��]�׽�2��$d�.r"�n��&1����"�
�8	�*�/�P�A��䞐��w=fY0�����VZ�4�R�F����p���q,�����m���gy�Lks���UYL��,�@��J9�FW,�c^��HR��O�,��dI����MW���M�{#]%P5
I�$�
�0";���ǿ���>�����RD98�|�e�Y]�F
�Kկ�jzi��Z�fI����� �}D<�*����g~<E"���\�����a��:D��W�������&b�|Q/��h�k-��0�ʧ yY0c��w�=n��+���w�= |��D��~�O	��:�����k��Оw4�+��i����|��-�$���A�W��V�$�X�.�P&aRcnD���2S�V�%ӄ�@�b9I��`�fG�����m�&��1�
%�q��򩤦�;\	�;��>{����/�����W�����IC�H��c�&�]8u��/r�s�����6�.��2������E��.i�.�kenO�_'ͳ�-�0����Qظ�[wJ:�$��ZQ�9.���̴�Ug�%���`�X���?�+X�fZ����"���!�ˁ�Z���_~a��쌅N�d��I��I
�@��tEU�a4�qayp�垹���oM��kÇ����D)�:�VyM�	�Z $|�`��`�!/�y���y�mJ���k��|`{�o�Z�2�_��x��^��������\�����ʙ{/h��(����5��F_�nJ���@nŖ��\ ;�d��NyV����7��9V�syr��YOY3�ݬb�\М�W����g1m�?����p�P�Do�`6�泙��k�a�t ,��,Dֻ�v�w z�>J�O�$�4��*�VNsPv��=�����|�=~}�B�m0>���X��m�e(2�?s�`�����WS�q��"$h#H����Է���c@I5fH1v䲸��! \�5�'I��q?�W��
v���up\V�Ƥy�}��J �VN�xz�bt��5�~�G�G�*�Mx(�,��,�
��g�_���A��
ٞ����v�pq������&M�,=�H��ub��˜[��Ѓ� �W�b��-��������c�gc����2��ov��P4�!��H���D`�R����3�>{Hco#١��)L�\B���KYnq��Dg�o&�!������+e7�3�gBёf�k�\Ⱥ�њ�+(���UZ�K�zh�[̼b�8���!�����;i$t�r��G?$���^\HoXTv5�O70�S��O�0'Ү�rd|�"h�µ�ꊼ�a>-sAv�I�T�uR�,��p��M��NC{rt�%l@(�^Us��Ej�p3��>���p�s����$,P	��[�=	�b
RѾ���l�*ӎ$܄]z�_5o�j=����b�`�Wυt�������~sxݦ�SJX�1S_�X�ޮ�Uwސ�#;7��5�+ݒ�6}����)�BdX��iBVVe�4��^b�{���ࡶ tI{T	f�lk9r�~ra:\�)��]*ň\4[��*>y�����HQ���.�������K���<Y"�Ea{Tç8��5���O��'�G�����R�֐�Y�_N��M��Qњo���d�����V���!}�����k� v�[���:�>ጥc0#�����l5t_�����npDJ\#v�7
�;�tv��c���O���z�Ӟ��#�@2�@�����^K=[A�^Y�Hw"�����w���82<ξ����^�qz���K���El��s��X�Jh�s:�j���%�:������lgے�p�Y�U`nc`��9�[� ��j��M�;�AK�&O`�K�&MU.j�-�<�yo:�P=w������,��?��_�7����3�ϗ���E�l��K6��]��2؋{p���;����7�'�=l���PȒ���!�Ku�z���:�&�F��Hy�:�J�=��I�	M�!$�{ĸZ�͞�:0�[�h���`)r�賕��U��`���u�#�KS���_֯��,?>[�r�n��"7���"�+����.�|��T$]���M�ӯ��
�FU(~��`�p�(��5�f{�|V7S�,��K�XݪQq�-��]��� ���N�챨���k<��a���XlxV16EB    fa00    19c0�g�
�!49N�2"�"�P]L�d����F�br{�;@� B/:t��H�bx�}/�_ �@������,d�.|�'���%A����E��w-����7g>7a�1Ϗ%`e��ȡ���5��q��*qa"!f�L�� �V,O�i.x���2̫>�ͫ<�a���{c�d}�Q�H�Ŵ.��rP� ���W���n�	��-|�^&m�Zb�����c�&��'-��\�F;�� R5Ԏ#��f�"+��1�:�3�T˕��p�e��v��5���̓N���A�k����
Z�P��V�_i[i���rq�[�
R��k5���i��@.��q��>�$�ҵ"�aӱ9K��݇X|� �M��!���xR����S���ZQ����}�˝���q�3π	��AV�
s
Ϣ�[(b�{o�ۦ���Y-�̿˚���
'c��x�լT�$����Y͕�v��}5�'&��_�W���˳u�����Sm�Z;���R��L��9j��7B�\�XQe,��v[◶��w��B	B�+�[D\Y��k�Q�е���-�{���R-��/�d���J�x�9t-��J2ύ:kZ��(������PR�'Du�d���tBZ��s�s;c�|u�roX��cO����Ds���)�n��r���R?�FW)�T�����ʾ�zN�F��Ȩ%�����O��S]c���ڭh9��^on'���'�e���\�ͻ;�V�YQ�}BMs� G1�ua
E�ѻ�)tI���[sj,�8`Cz`Ҝ�>p��Q6g1��2�=D�T���|{*_H���ڏϾ�CGl�gB3��;}���d/܏�@=[�βu�{�I��r����yJ�!1�kj��ܰb�~C�����g�-����ȶC�Jt����N�M���5���~6Ǉ���)c��u�ט�3�S��,��Vu�㜟��U��v�6+�Z�Gm\��R_�:��@�#b��v!���.RIL��ND����&y}ϴ@��]��XG�)�0��$+BwMA�]�1�{Et_�,����F��ةI;� ����K�OI���I�6���,��糜n���ˮhiY���ȉI׎aK�Қ��0�Y�a� �Uk�}9���"�;�}��&I
"����Fl]:@&$��/��a��;�]��+���o��z��Wܞ��bC��o���~p�
�_^ Ss�r4k�%��g��&Z"��S�3�"�Y�$�Ty�X�0��5���>�b3��a�T��/���U�U~���i�/m�s����t��D�w�c�Iό��r{]�d��5^DU)���\g�[]�`�i��z˛��ܺ-	�9�qw�.��ض1���;u֏̤�S��!6���Pg���U1!����ox�|���p�9�����j}kVx�}o�%MijA����c�uxi?�����g��3\H���J�M|���IG�1`�cR�_}���]���=q z|&��w������Ý��a�.�I�ԕO����L��2K\���i��6��&�'k�Y�2�Ѽ@�b#�I�� ���Ҥ*��f��J0�
@�;pKo1��{�	�����`�w:WLPk�({�/��#wϗj���H�a�_�!�n�c!��:`�	1~	��N��5�|�wn�����aL�����+(�.��e�C�'�z��{o7[�',�O�T]nnͦ�Jn��~��!�,#T�=��hp��U���8�]���f�/މ��W<�z���c��n���M�D]lYU�t*�G:��:�_�]���n�-|��҈���0u��^%v�"�!��`��T)�25�nx�T�x�(w�!�t�,��l��p�U�����ر�<)����\P�j�Pt��F�O0�V��K���޾V��Č,}A8*�2� VR7��7�a��M�='.Nԇ���%��K��� .�V#�����9�y���??�/�?"|.���U�A�h�⨬ǆ?�C�=v6}�Q>��%A���g�n!B��a��@ Ă>5����-���ߤ�h4���T ]�a��j����OR���ɵطg̢��7�,��6-��⹬Z��p���j�����U����a��=j����Bl3t�B��G�Ի��v<�c��S�wޞ�[�,G��Z�=x��ͧ�����/�.RY,�g��eSv�L_קD��.רoPD������'�6Ę_���z�>��-̜K�x��W ���#ү�L?��VC�	I¡�([���I�|��h�SC1ٛn2`g����Y2a�$�楡�<|�CU6o
5�9�^�*N����f&䇌���z��oD�j�ëK3�lM��麴�ï�  ��8��0�=W�-�t�nM��N�GƦ"�ק��ׄb�	q��2�?֚���f�P�s����i0��M 2\��zʢNÂ��V<鞟gL�S캉Zc�Z"���b�z���[gcȻ ���.S��\��$m����x�jQ�A�:|�֓����5V�J�=�HW2ﻱ��J�_4��
�)��D�_)���"�['/<vAg�z"#�}w�zepUpto�``��
	��;�7p��K_� ��RA��˦l�c3m�U=\Xǩ�p�Q讼����7�{��, �/�h���BBkȝi��]5���[��Ng7akj����튄~8[�ZE8,��U˹
s�:���S�U(ۗ���z<��n�7si�}6W��f�{'-j^�cǸ	D)K��C�Tpo�"�)t�?}���@��YY��~ˋ�yl��_&a�� ضA���!V���V삌(Qh�Ӡ�P���=��J���
�e9>��O��2)0��f2���v��5p]�y�ՠI()l�`0���Ȇ�Q�k�2��ɥ�F�v�6c�/�Ɯج�vs��R�u?zǿӼ�pJ� p\�Ԑ��-�JkTT}���*��s�V����vm#�6��I=�Q���39N�t��sև��A�FD4s`|���N��m���9?�h�y�����8��ϧ��J�F㝛����q��=���ƦDhM���N��
5��H r��2	��r֋̃��b!	��L*�cB���a��J�H��}J���-���2�PtF�p�XP
*��Ww$�*�`%�ض�j:�h9�}e�'��Sͤ�2�΁O9���^e��U�O���Qq}TN{�@��n��<7nT��r=�)���سl�t����2.#�W���}TQ20�h淼�u�o�g��%���cd�z{���;i]x?�7hs�U����;�% ��R��d�[ΩڰM¬���B�R����Su~PxL����j�*
oܨ3$'> ֻ��E5�Ɋ@���^��<��@on$Fp�&
o�pPr�B�f0D���X��M�E&g�=�n��-
���H{�߲l�;���y{N��
��b��|Ԗ6�����-N���I5��b2�=ݻю���&ʉ�XWF�o7�!��>z-zB���̫�Y��l'�N�,F9�r=:����,���c?�a!z>G�XB�Rw�[qgl�&��x��i�����p�@��h�*���.tA�a���4W�kB�a*�b�Z����Dfr��h� Z$�=��k�%����ǡ��lt-�XEu>���� !��ĝ9�F������-�ڬ�#�P���W�A���Pw�J2���3��7Ӹ�K@�N�O��'w�7�e��-�� -�bJ�|��I�:|��HC2�*���y^Y�����������<t:@��B�|Ķq��N�DN����q�7o�ۂ���je�?t����B���9��Gk�b����. ��x���
��B�$-'3��z����9��dz<M���)Jv���{NMi�y���@�6�?B�^cT�#���Yz_��;)n2�R!rI�C�+����R����AP&!ٍ;L�.ty�(�/�X�v�zI�.`U���_�-�-wcR>aI�o�������gI
��+L	A�s�A�n�]`;i��� ��0��h���-�V�)�+mxL�O�bX$=ZAz/5]��u�ٯ�H����K�$�	��K�cgHgW���)�u�|���l����&l�z�)��\r�%�����4���.�+H��Z��w��C��������ò���\��F�B��?6|�
c��Fo�P���3���ZV$�����Fr��pǴJ���)����|��:������uC!�,��J�A��S��_K��q=`��Ѭ�"^��|����v�J20N���*���fx�����#�R��ۊ�	*z��Rq���Tx�א"Fk�65����.�S���r���韭%�F��cW��@�-Q�*/H7OFb����<��'a35�:-��q���d#�}���w��A��B��;�Y9���Cu*J���[�@�|�E��M	��W�X	2ʽ}��������3Ho�F���t�7ۜ��ʡZVH�V>�s�"���lߪ�-�8�b^(��$y�l�T	��=���q7׽�����mq?���-*�9��-2M|��3d_D9�g�@)qoY���-��m��z�������i�%��Q�F�����O�.M`��I��h�5v�/0���ٍ�����[�<ERܥ�T6Q}��rҭ0�i�P���í�}��U�'�������r�Hs��P!�MhΆ]րj��9�H ����$�������˹�aU���|�J���<��M�"U_�wk�zR$�2P̪@�S�̿����F�V�r��=`�*�1Z�������~0�g=a�D�Z<�Ǐ��){�O8�,����Á�a��C?��d�����t�;w;�׆`�id݈͹N��G�V9����4S�	����g�д��SyB气?C}<>8�'�g
�o=��$���J{�qM�/N^Hf̥lPE�����5���U����Λ�>��C���(��\|��{���D��?3��/�� �2����=KQ�r��*Ō*`�e���R��y����k����QP�[	�Į�2ծM��i��z�n��k���qVN�O(���7(�Rn>)�!c�p�'W��E�Ԏ[�!�|FZ����p_v�x<+GHw��x;���M"kR�;ԗ{P��<�}49²�֥�p>6��J�
 c�k% Y	(���X�8exE���Mb�NU�`��4d[�*R&��Tƌ3C��O]V��ɡ����'2"��	Jl,>�l`K�V�ʞ0x�X�8ò��%#7�[�<S�M"9O\(_��١��H���(6�s��s��8�����/�1�$��N��t�h�
�Gd*�΀*E��r �1 Ω�VN�w�Bӛlu~کEl%R�AwU�n6y�zh�7�B�Qq�A��H9
�O��^#����~��ͩ�a�-����[�Xo�� =�tS��@%6H���ŝp'���8xEi�s���5�([V9����ew���k�v��*�k�{���XEu�8j#�w�ᑖ����8�ϰ-��Ɲ=ܬ?�.�!�6�hO����2Խ���E!�ب�~𠡗z�re� [�\x��A���~��r(6}����W?��W(Ty�y���H'@6�d��p�����ni���V�X�EW';�z%Hg$��b���R�P�^�������U����o�@w[Wl�Z�H?��c�������<��
��C:�m%�o;�c��YP|��/��vf%暫��i�Wm"�K�+I�Zm�����!�5�F ��ڞ]Ȫ��Bs��~��R�þ�^&_�K��]=?��b�Dw�./��zx{��Ƃ��Q�i$���8u��Z����4U�/�g���m���F~]x3�2�G�.+R+F�.�aTA�e�������i���P`�"���F`�hKK��b`��K�>a��ThH�p�L<��m���Z�Jl��a	���I�:	�8���I��뼕Y��>����&�6	Y�w��)����|��aD��hפ�z�T�Ȏ�Цt�[�G<}_���s<��9�=�E�%fj^��((����1�n$�>�T��yz(��Ŭ�b��ߤ�eu@!J#)	r����v*�N*��y��*$���3���c��K mDr��ŭ;jj�!�=R+�	��B	#���_ Hۭ˓wԂ�F}m X���r.���3�EX/��k���9 �G=������TD����p��W�Bb��`���n���3J4�\����p=��]�J�u�*Č�iκ���A�}}O1�&`�m-�,���-��k44Z�%_L�����=�>�^���:��U�3y����oD$���m+����P�D�i��0��t� ��C[m�K��U�I��tre{�W*T�c/��jx�+��)ɡM��|y~�Ku�^�7�5Wd�x����%��9�8#x����B�ԋ���v�&�=Ӏ�!R�9��-t�l���B���Ϝc�ْ�Z�N��@��c_
z����XlxV16EB    fa00    1680�����$D���(�����c�z�~-�E�)��l�:����Zb6�ê����7p�X�����>�(�&���e��p��W��C�j{�	F���J^��a�|�#^Z�v[>�f��� ����]���p�W�8&W}v�:��>O%��vY%a���;j��%a����je;�J?�@��FBka%���*�~�l�%�Yo/q%��<���Ej�CFҧ=���V�3�yM[c�����N�~g���@�oJ���r�:���{�����}&�w?��:��ޥ�+`�m�� iH�2	SXs����ad_t����U��|]��V�8%G��إ`8 �ClO��)&i�z�h/��
s�P+���� R�J�rPbp|p����ʜ��O���i	���ٓRb=��sZ���-��#c�	V���Z��Ρ����,�p���6��E
5Zqӿ�,[M'o���4$�����I�9�b��9s�ĺ���/��V�'j7,�>���Ւ[
N�CU���Y7�Ҹ,�����X�K��[d�u^O����>OQU)�t�,1q��:� ��"~������i�|��y8zj�L��]��ً~w�Ah����8�{��_���ٻ x�=^Z��'[�V�aŏ��U�l�p��0����y��dF�o��|�d� �G��@AMMSh�Ά��h�0�u��M��®��(���j�E��d~��q#�х��Q����k��w�M�%?[S�5(S�����f9]�
? ���C�XDO6�Vn�ضa$��I0���>j�MmB�����/����cV	Ws�)Y��J���䐗gX�����>q�)9\�nJ�5tD^���	.�;la���xø����boht�֪����o���󑄃���l�� z�ve�n�ޠ��6�5<�+2[0��z��:\W�%<
�6�x��u�RLx�051��5�3���: �(����"*��mw��G�7� ��`AT�����d�Xc�����1������3�E�xZ�M
o�`�r�7P�=b�/Âi F� �z0ҝ��#�8=�;?�u~�p���T��-�>�`� �V�R��Qv@��:q4MGxY�( ��<޷Z%�� ����#n��L p^�mY���
)_����X�ʶ+�h������R��f�+sp�W����gQ!�9_��J�6~qțV6��&��;�2""	��rPw��?C`�r��,IOg�R�/��MM.���-��8/������r�#?��g�%��m��"*�96 �{2�%J����s��9�$��d쪺P��?2��a���X�� �3�p�`:�k
�(U�z!���ea��ZQ�9|����S�\�*T��b�9�j�`�z||��6[i�N����g��湽m��]~?��0�����^�G1���$YڍLf���@��n�߫�7X��r5$�}�[�'�*�(Z��N$�����L��n��m���F��:�S��!�KW�c
X����?p�f`�e��Y�x�a���T�A�{ʼ������AP��R�0�{y%g5����+1�Qcq:�4����'*�3���E���h8<1�������2��P/}�m��.���&�:�2x�9v t��L���a��b[����P'ĝT��e�pk��W��z�5S%p0uuAD)ys�a���C�NH��'��b�
!�y4�8$�K���Ug+;gCp8`�@�m�Wi(��������1���Hee�n�y�|���1�����Wbx��O�0����&�
g�����LɯI�A��l��ۢ� ��]z�?�@�����G�(��o������%�a$Ļ��YU]5l��AΫ��-h���ǫ]�9?�P�H�����X�}P���7ҥ���o��D�IӉ".�M2\������&��>�j����{M�_`�o�8dė�[��PC��ސ#g�p$��]K�/Ϊ��?)��w�g[U�bq����И4�b��O�?h�l;��9�cw�M���W:��kTVWV�1ر��xzE�F������s*��nQ�!�X�a�դ���p�:��^b����s��R�$�׽�y��3��l��/��C���إ3S
B�|C;W�!7�5�,�Si>��[V��Q~�勲1���n}2u���:$n����M��X��-�34k��r�
�T��'���V,~gt�ٽ�?,�
Y��c��ص7�H�>�P����(�OF��B��D����z�"�*ۈ5�8W	l�>d�/s����_�ʖ��U�E�(c����6���B���W)�Wj�؜�� =��GX4�I��\�*�>}�[�6o�C��ېI׽QbS�"Ż3Y��ڥ�ߡ͙;�O����O�$�s:G8�I������"l�.t�{8*��J6F��/z�nD�ɦ���Sƒe�����W�"E�����j��@P>q�"��������.
dEw��S��+���r���P�j9p^@
���70��z>-�ӂjX�.y�a���~ַ�ʬ�||}o4�v�U&Ss/�<F��L	�/q�v<�Е��i�E�bT�`�����A�֡[<��z�L�--T-� ��a;��GEW� a�k�9aCfw<����D��b�_ʷ�~V��$!V��O.c�1�����8�G����Ak��{�9=L�:>Z��s6s�� .xM��� ����Оv�o�08�u�l	�ޢ�G��Zˠq_�e����OjE%3y��bC�`��\s��%��<�}ex��TƷԞ��gE���3�4}��WT���gZ��/��?��I��*^��ؚ�Q�'���`�.�^_��2G�D��Ď�%ü^��v�>�����Q��?xW�'��v����6�㭵W�1q���Az�:?��M#�-��|�Z��O6�t��Ph��̳}�W��R�2��GŢ�����k�|w�?�d��r�z[G C�@���辀@n��sQ}�]��18xx)��H@R�?QS��}��?�=d'����9����'����~���6ly_m�E�]O�����l�9"/�T�!3���x;����3βC֙*�����TZr�Ҧ<뤹d�2�+ry�BTi����XYf.�r�,�������^�_؞�ީ��C������������~��Nd���<5���0�j6���5��Q���G��)�fJ���(*����P�y���Z}J(f�bO�I�5Q�КS���*`]��&w=�B�O�ߢ��u�6r<��A�0s<��	��6gq3K��k����P�'3|��7�Db),~��Ü�"�I�dr�|�~��V�$ܜJ���D�m#%��y[�*�B��@(����ETYzJ۴��n�]S��Q�Ȍ;@W._��\�����j[�����Nr���c�5#�O��b���u�� �z�^�X�7`�!�����_	M�DS}ٻ�Fm�=�6Rf>�A&6g0�8�8p�r)�
��RX,z����V���;e+Q
T*c��N�X:��e󨌒���v��Gs~8��a&���X`>F^0Q�#rG%�KHޔ4<;��uq�?��}��ȑ�*b����v��6b�H�Ő��=�z� {k�t� ��*�x�Y�o$v�y�:<��X9����i�$m��9��YW�X�iE���1�8G��/���_{ƺ���c�ċ[��'h��	(���sFT4u�8�-P����n�!ĥ��t��`���ù�&S�;:���Pt��8XVs�?���eכ�?����=��8L�����-���2oц�,ۗ�[���O�x���`8}Q�y���h:C&����Wy%��=�����,̀J/B��hU��E�1	���iHV�؇w�{\�}���t �N+�� ��я�y�~&Ћ���cU�.���tH���rEۙ��z�9!�8�I͓b�|�ƐG���D8���-2�<�ٴ��E>x��?�_6�UT�ʑ�9�C�&�F�V�k�AM{,�}o6<f�>@�6�&I��rUx���b������A����55	�V�v�)IT��o���N?��XIPN`^���������w��b�6<����D����3�Pl5��;K���e�tH��(�������6��o�C5�IL�԰�Fcп^�0��,�O+.���� ͘+�<&w#}��h��T8�j3�A��鎰G�
j�Av�U��ד��h�3E9+"�!�ogWP%ǻM6�����\*T���*�s[fl�p�l)�����Ȼ�������	�f)[CN�\��;3|��*h^�M�3ꗼ����90�?��VΗ�*����m%cth�%X��&~ݽ�h�ѝ]F��z�&&�e�@S 7x�<�F�J�R�./�C��}m�}��N����8lV����QP�\i?�$����{O�5�!��E�*�=� tE���`Gb�z���6o�
����(Vd���5��i���d,�Z����C�V�ͯM�ᾼ�CZ+v��B�񕰭��K:�&��D'.D5�^Y��q��@	^2��Yy�o6�~�te]�˝����Q`�IŇ�e���ű�o��1A+�O�t�֠Y;i�Y6�êBZ�X4n����]6�>���ѳ�������;�pS<đp�E\i���޻#���'a&����yv�fqwG�ꯛ/�����Y�s��M�<��>��N�$�k#��bƘ�*��u0��-�sQ�aےt��Vh;�.�Pm��#� jI#���U%>z���� |���iZ�e��R�ֹ�A�0�w�Pm�g���ڤ������yi���"�4j+�1�;�U`�!�9�Vs�3��:`���9�S��3���i aX��/ߖ�b�O��r��T�@����:A� ��"y�g�k��W� �wl�5 �>Á4�uA*�3�G�|hd��]��왟wP�:��07��
a��������г!�),�dY�د�I��8�:a�&�7��PܸmhX�b|��3������n �5�u�4d���}�3��d�໔��Ӝ"�o�8֭�������|i�mFc�c��ś-�f�J�p�Rq��v��!Q�;s�<�F!�8ژ[�8�X$�TЅ�4h���F�'0+ ���*I�u3��C0a+51��5[��c~�D��	��r��3�O2��a-@pg�1Y�<��Lk-�fֹ��rWM�����T��U��~�!?d�u!�2h	�ed�b�a��]�[i��)ʯ�=#��eT)�r1��ꜻ-'S��]����~�xc�Q�2��Q�m	�Dͤ@G	q(�*`���>��yU����x\*��V�������Z���@��1@!d���&�Ͼ���$,�(z��+U�gF`�d�1�?���B�<��9Vv��S;_.���Y=���S=��Ba��,�cxm�@ ��&+�(��H��V�+��� �]��Op��1�<�����l^ }�G9���G��#�K��D?��Z� ��ꢖP�y|L���ܨPI3�O ��gYQ�����k����#`��p�w�����I|���2�?�]��Us��~�e�����6Ay䱰�]Ê�f� �[`6B��"lqN�a��m�%
��n��>��5 |������hk0g���WY8gb#��Ϣ�� �΋�m��J6�3�xO���:t�+�ܭ:OiL|���C�=\@��\XlxV16EB    fa00     c40�����o/G,���v/%�c����z�!�?�����ԙ�6�ZC�����v,rx���%������P�#��`�qdK��F��DO�\�<Ѽ��p��D%L�␄�>��,��H�Y�?��9=�L�����wp.
���� ������ihr�����x�SB�*��֟����䵑�u��]q�Q??�8{��!V�{Q]��n���ówY;i�Xs�R��z�F�d�Ȅ8�T�g�x�; i� ��GЯn�<خ~��S�5�vFY��$z�e�v~��F����v�d�9�3J���-�~���~ټ��0!|����ө��IU�N��ߍ�>�C)��6N��g�B=w����[mCY��ڍ���'z�RwD�2�E}���n�9u$mժ�}h���G�3����6�D��kd�9ĿDÿ�:Ѥ�:Bn]��5��E��xƷ�v��W9�ߟ�F�ؾ�w�{!���L���n��9?w��=�;Z;&�ei�6j�i^� ��i�[�5���Q��*?2C��&�\���ȍ���XCb�b���5�il�N��2�h�ԕ��lB}��%�w9Ϫd�{ \򍃃1��E��MK���[��A| ተۮ1b�F�BU����Y&������@��p�N��X�F�"T���~@*��)l����p8x\��F�D�mWfq��3�
�_}/�.)g��*��,}�:
k��b��6ɖ^���~�
2\��|GFU��Y�䋥�WEPPK��Z�}m�ܜ�?��#����Ȗy���*9��'�CΥ�m~Jj��X��c1�8��  �È�*H�I�h��D���G,����P6w񄉵��
'�¥�����.�����I{L(ޢ*�����E��֕��C<�h!��n�R(����2��&��l�k�	���㲼��k���/>�<���
#A�����\0�~?�O���_�Hw}��LC�Ti?4�~_w��1/ˤf%�I����U٭��Q�7;s���Zon�i���w��c��,���m
(z�jE3^kQu�b|��W�*���x�!"����k� �k�;xj����Tp�M�Z�����s2��v�Z�U������䮐�z�So�T��~7�fT�t�� �@1l�'�-�T-���'*��Eok/�m,C��ƾN�o�;����4؆4�קn�K[�����6}� t��̂����B4@[
��Jl�,�Jiy# [R���cӅԫkYk7�c����-�s�pc�fr�6M�n�>"���r��@U�,�="weOI�f*� �A��GF�A�η���9��_v���R̅�0��	�Z��+���:ߘF4� �l��X�+�~�q��g.:zx��MX���@C�P9��@���A.��vX��YS��R�K$���4)��݀V{�:��	��i!��;�FH�<�i�U86�3����=\�d ��k߱�S�6��ٵɀ�?	�����ƒ�k��6 ��x�m6�Z58���^�p��E[�v���xb����
Ԅ���o�ݪ}�\u�y��9��;�Dדj�t�d�YSS�a��!���۳-���-�v�"��Xd��e�\[�n;"e��{�>����&wɉ�t)�S�)���>�q�N��[�k�,�V�����tO�c����̞&��������aO����4Qh�1kAq�ۅ�z����q$���eZ�-�J}a�rr��O�ײ'�&��쮟8;�p���)�a��-,��%�G?]��G|ަp�?��}O�3#��B��Œ�G�s�@�P�6L����oeO����Ɗ�z�*u1d�%}�z�8=|{�Qd�B��`����R��-��Fr�H�������YU9=�B�nxZj���:|�Ơj����S�`,�_��o�`i�ل��R��b#N���a6э6��e�e�wx�Ǥ�oT��԰�iAJ�|��ѷ^��)$�$u� ���h�"�$���i���-^3�s�a�)c�6���|w��*�����Ǳ�aC^���6s_�x�y!��"tǽ��J!��Wݡj��gl��~�DJM[�_s�{h��ӹ�����Yxa �B��3P�J��<7��6�Y�w<��9��<���L�[z�O�ѳ*�T+� K�?�~C�5^6�<H�y�NΕ���I�:�ѳ����5�BX��w<���P\(-"\�nR$W*�vF�~l`!���]��%� ��Ƣ9WS�Y��`/k�$N+[��x' B�	A<��m��	]P���������M��b�'�w�gfZZW3�*�Ÿ��[�Xˏ❌t^k�z�KX5`1�!��8}��}:����Y�pr@N��&`@�����]����8#�;ຼC^[����|��W�HFG�<��=t�ي�ع�t3��V񉄣_�1_����w��Q�%�� b��c��H�(,�가4��lc�����~������ÎY���c�mh(a-;��ƞ�$��e�4_���G����\����%�h�
����=T��e���8!P�_M��	@��:rш��d�e�*��"ն|~��O�jR��6��?�f���e�)��첑&��}��'��ю��b
����s��?=%�����!�]��;�Z�p�u�IQ���Gw=����?�X�2Sb8hC�j��b��&<2Le
�DD�H�1�%���8|ZC��0��0^�U��1���;}�� 7�b!i�e;�P�rH�u�]�J��օXTk�ߨ��I������NN�bJ���Z�#�Hp��������d�h;�!���.�q��B��P�5Id�b;�%�h���W���!)��?W5���������6�;�gb�M.c�x�/^զB:�5��fZ�@����W`�$�F�=��w�KF{J����,�g�ܣ�������Ȩ+���M�#���.��yB�@�ݝ3^�)���nĵ�U0�r\�)"��k�C��˶0D���b��}k�����R|��ğ�@�O�#�Tcn�s�ܖ:&�@�.�v���N�Gn�5ı��E�W\%UE�T��XlxV16EB    fa00     650HKzp�����R�S;^e������"�^Qx0��|%n�^Wuh��&,��1_-��4A���5��JCy0�3�n��4S�1��V�v}��8��C(?C��u�ƥ���;u�����T,!l�5?Wױ���Tg��ty|���D�$w����c��'��T���n�#;�٧�_�3�s��"B��pn����Q�����q��e��]�7��}�U��J�v�1�����F�D@�����!SC�8E��U�.Q���>T�i�9�@��2v��X^xZ1�AJ`^�L#Zd���S�`�W?�dRv��)��4�A��@��̷s�^�0��qW��y؋d����E
�Ù'#Ɖ��w
_�1G�k<��~�N������`b��|�{�E��f�\�1�Ϯ�;�Qg��$�o_}��;Ҿ�bCF��~��Fb�/=��$���?�/ߞƛu�0]by�{ �:3�c������9�4��p���Y������4СP�a!%�g�hiF���4�5�3���3>�3�U1�����j	WO*��Bt��o�;�4�]�_�͟��FVo߅m�K���	��]��WM�.#�-��q/��B���"��ˉ��H�bkA_��&�����ƆPa�ӥ�L��\�1b7�Q{�f�t�@٧��[j���L�Ds�s������0�[�<&��k�P�7~\������e�H�?.�Z��,�oi>��>�<�p�	�$`����q������w��峏cBL���*�����X��¸���*��Zx[��5�/�r�?P?��,mD	��ر�)n��hPX�P���x͡�a~��Qz�Ȉ��M\;Ǔ�v�d�IJ�i)�&x�ѼƩ��ǭ�*B�k�Uu�?��V�_�<1��\���l� )��%LG!�k<�J��F�$��=3�=0�0XQב��� n��b�U�駘~�p?^����}��𹲏�'�ة�x���Tɋݘ� g�;#��S��aa:t�,N�$�_]�x���r(fѭ�9�Ǘ����m�TV�>b��'�<ʘ+WCa�+=����� �1oep�I�ǳـ�7O���˓�S��9dq
���A�7�Ш/bq#�'�$��ս�d���J#f2�j7�Ӆylý������������>� u2q���/sp̲��x�6p�|�6�j���pl���>Qx�/��2II�u��ߪ)����mc�l�\9	ޠ�|�%����ґJU���Y�w����p�"���{�_W���e���Q���U:v�d-X�m��J���o@����ۄ�p�>C��Vcܟ�&(�X\q
��8C�#��h+�UBJ��O�u��'�'R��B5�z�s-�ml#r�)�4���x������kЊ���G��������Ci��\�n%�����|X��Ȅ���X_˟8Z@a�:��ۺ!!g7�2���~`4����o�o9��{v�MY�1kV
+$r����أ?�x=i�%b���o���9�����i�� 1�<�B��I�n�/ϳ�t,�t8�N��<c����󖠷o|��t�w$�s��s^YOM���]�a#�y�6^r7����XlxV16EB    fa00     5d0H�&-�ft~��01*��\;]�<�����H@��7�~n1>�c/���e�=XK�}�5sq���<91���6�	���X�Z'Bwy��߈���tk�ӏ�3��g��������Yf�h�����OZ�]o��Y�
�؏�$��$~n��o�~�~�=� _�^�h,Q�*\����T�O�a�����|���z��G���7�S�$m������循)�j��9�u:��1�h�zv}r7�[�r��p��� ɮ
^T�����N#D&�G�^]�_��>Ֆ�S�m1��ғ��O*��+	vS�X��i�5��g�R�m��;,�2����Ӣ-Wx�*�P�N6�� co������2��z�Jf2����0��v$� 4���ePY�@�@lr4h�ǫ��{�F�tD�����k"� H)��p�z�Q�Wh�n�g��x��x�(�����撵x�o�m���0���~��X���$[w|(j64S�nb�������]��Q�M��΅`	c�I{g�Gk}	��3 UQUw7�e��5��\@u��	_�l���[}$��T��L�Ak :�]�y!�?_Iq}�����H�t��gm��!sh5#�7�wX���9�A��F#m��.�#gW�?¾�K�
�v�n��l�$=�Dn4�_E�,i��;���䩸����Z�������(.� )WLן!/ȑ��s�����ꪙ�Ě ��H���j2����[�;��r܁���$	�����ņ������Nw3�e�G�P򖬽�c�5)��>�鑫h�9�t�7ۓ@�ݑB� BZGU�_���FSNs'�
t�L�<o�mR����o��.�d]k�V�E���@������0�����ʗ7��/�� (�c���/p�b�)�r:����w���J��f_��X�,
	�#P���إ�<*�������@/ۓ�+&��}(b��y��ׅ�I<�{j��� �У��k�Q
 y_�D�u�bC��)W>WyYY������-���M� ^��|@��zw���A%�P\0��J���صE��ߊ��I���	x�]��"B.	pʙzd}۳1H&����z~03ϭ�L�'lW�ġ�+V�3Kh �7��gH1uDX�IRN�<���t>ݗl5�tO � *M-'��~#C�{����SMWFv!,	��V矰�m�,F�`t���P%�2�����P��5���ИՆJD��m�-5���p����Y�\+��8��}9����R u���bf�/�WS1���_�xe�/d<��)����0E[��p&��5��QXG�'/a������Z��6
��ߡrou��8>��mX �/�o�x�g1sbu�;�1�3�^��B��D����|/]zB��v�3��Z��V�X��C떩�5�[@ڀf3VsM-#��߉�d*2��a�S�~�8|�6�Q!�BeɈ�'�����,�XlxV16EB    fa00     5f0@�`�n3�b�ݳ��#�ts'v�����U k�*�|��9��_/ԗ7��䐰�t��9��gt�lh��3B9έ���9t���t���Ƨ�K]�4���,���9&��^*I�j�љ�����'� �k&zHS�:/߽�8"O���{���u@�mf�kOj0�2(�:HD��^�M�׼�.�PW�r�"g��ӕh�h��� Ɖ�7��O�l×��qS烾F�ӛ�)i�&N�O��7�<I��`�7�<�t/�ڵ��g�B/n����V�lMţ�j|w��Ώջ�neD�Ǝ�U*s��ͪ��WŨ��
�]��-L��IK^.�����e��n�Y�b �{�y�;?ߛ�n_��wQ��	�iU���t ��ڪ�*f��"��{�U����R��O;`��F�"�Y�=`�
� ��Fi�|R����L�{j�g�9K%���/��A+~����]J<?��i�Hy�{[(I��#��g���t���P��}ݾ^l^�Ŧ
-���K��i�)0����b;vU���s1�@#3�xս��:�wY^��a>E�(�,U�L�9�� <�.
28���B/X_g`�rYyQ�8�Q������kt��:�hӆ�4��.�BF2���S�\{^af)�ϱtl�k�G^�S�V���LhC|Sa�O�z�x�b52�HD%��|���/���ZĮ�6�����KP1��>��1�{f�T�8�A����ިlw�γ�^-4m���}e����M`�}��ԅ�(��j���RW��סt�/A���f�E�ޏ~o<|x�ص(��r�e�x���J�E�i}�)��_+�kJ��JB��:�5&4v��[�rp73�˕aRO[�JX�hMx��܃#��;'T��8c'o�0~�*�L�+8�Q,���x4w�V�;���:�Um�"6��ڻ�V� �S��߫�[��%�A��ϰ*U��'E|T윧�ժ5�������Yl˕����;ܪ^K���_ǲ�_�G�n8��QaX�`�q��x����<J��d'��4��R�d�d��HX'W�����r�e+�P�gx��Z��E��<���ׅv����%���)��\%�k.Y�c�~�*�_"&p���7 �fS,('�}��s��0y�yw`S�+6�*Q7�K~3!�>X�"�ܕӐ�<�CULB�b���� ,B��R��C�0\�e�/x^���{H��+n��7�#3^\�����/_�C� �,�`�vN~}'E"�3�	,�67���6�'� ���&�i�W�{,����m �S��6x�9�$�&�[��T�_��2�GX�n·��R�(��Y�Qh���Mێ~DG�G5�]�o=C�d}�+)�6�A�h�9�̑>&�S&;_�V�TӬo�VǤ[�}�	�`��VȬB�~����z�h�, Ȉ֡%ez1Qb�~�������1��4Q�_��{�^p<[�yM������r�E 7�U��bm���]�{��V�XXlxV16EB    fa00     640�&��T�pw�E'���R�v�>un=H�����
���>i)��x5��ަ�i�h�~pFiw��yHg�EHNqJ\���ƴ����b�uծ��[���8�������i��Ե����>09��Ժ�뿃�p�Ia[~D���E�l���Ush���^���`��(�;9��h��n�a��Jx<
c.+>��$݊����ю�ҹa�
@z) |�zCdlƯ��ɿ��G��-_��]����#��R�y$�k �4���ґ	��5��T�^�t��xa�1>q�oÜ�����մ��q?+�.p@�e%A:A�B�mLćo��×ʘJ(����Lg���6��Ou�y��I�t��O�8���'m��"8u���m<cZ�9u:�G���Qx�3ݗ\҅&ר����G:��G�de0��҈ھG�<Y����]\���-D'�򘿆p��Ͽ���@3� s�$��
����V��R;�$�lA��xrxL��LA�ǥ�RĵC��m돸"�7<��~�5F;w��^���_���j�B%��7�w�7�4fG���
Lt=�I/e��Q��L"�ie�(��4�c�^�sb�o�N�M��#]>n�$�+����h�p�*��.!��BǆȲ�@�5��_n�/jg
�i�D�����.��w�V�ރ������K˺��\��أ �P=b��t�_R�kNZ2|��d{'�^OJ�*��O^��|�3zl�;��Z�M���7�o�K檐00��h
�����N>G���b�ح��R8�c���=ʞ:,)�b��A��'4&��K0'��*�q�rvC�_2����|����'n�����@�o���gE��6�/�~U~j^�X�Nۗ��eJ��K��{/����?:w ��$�CD�K�@� C_��u��wE�Na���+>��K	e��}cT��rNn�s��Mkf�2ū�f�������](�1��;jp����Pa��c3N����Z\��qV��VV[T;��o*ٜ�%M윢��"V��.ю��niQ���PR�Tۑ��Fg9� ��6.��"qlp�l��e�~��|�K;�n�9+�*L���tx��>���T{�L?&�vO���u��r~���7*9�	�w��N~p�K���gY�}_�挩�wx`��>�o^g������Z���pVyX:�����(�/{X�m�+�
4����x5�#t�\We]0b��K�'��01)f���oo*g����i�I!2�oNrB=S���������@eB׆Ҫ8�)�k�e��]7<��7�詍�n:R���k'�G��O	�+��:��JQ�s6z�$#����ޝ�h��-���`�e��F��j��&��j��!����)0��}��q��NH~b�#�܏2u��SK���׿�}��Ui>W�k�����E�{6�*�
5r���8Ik�F`W� v#| �����;и��q�j�P��u�`[t)�]�(3�:���G��P'������*�K
b�U��VU'��{�m�>Eѧ��w�"�۟��~"�i���8fs�؛XlxV16EB    fa00     9f0)1��&l�CG4q�'��V���4�,��1����,�o����Q*���j�S�A7���WZa�M��g������L'pA�1��P;;�����~n���*nvᥑu�m��F��5lG`(PFJ���v���ϲ�Ӊ1�0(}� o�y	���_>G<\����&�����o&6+D�[�͵oC���d�	^ŝ?.��V�+1����K�t.g�Q6ֵ$n��:v��0f�(��5������ob��0��Y1s�����2(v:�H��sm��@��Fv �D��ԋE#�8#��~�<�5�7I4ܖ*�n]��L;� 	Vl�AD�K;�G�'Ψ�n�W��i���(9t�h���^�Ʋ����d�\��ͤ��i�m�^�/�z!��U�"HNH8d����g��RwY'hJ�����R�!�7�m
��!h=��Yl˛�s��F�`	M�gusėZ��a�3dH|��xZ���ŧ ��n��	ǳ���(�gB�!���;�r4��&3����k�P r}�k0ȹ0��Sb�e���=�`�?�~
  �]q�}|��v/�f4n���1�Ƃf�p�Z�|��i�jE?{�$��U��NB���-��㫩8���}صё�D~�tř^�w��Q��f�!!�՝�}�GU/z�ezr�n�=���ᘭ�����®��.+�~�[��5��:��A�7[b����*�ƸЈl��ђAkֈ�c�����I���8���n�G�������'^���z3�E#�g�g�!��O�I���FԨV�i^�^X�Uz��9s�7W�q�qx�u�sj��8p5�ާ��~}�8�O�6Vl����o=:|��M>�����f�
�l�����*ݍ^�P�� ǵ~T$��|��[l��vE����߇��w*9�̲�=�E� �Ίi�.4�(x�u_��Ҹ]�� ?!:�B�p^��
�Y~�cZ���>�J�+����L:�$/�d�_�y�>xe;��)�J�����dtK�?�s��W͔̠`�S ��n���4枚%�$�D�K	��pIz��7�8�k_)V�#ކ2���{(��1d qq�n
�ht��u��$	�5�hɦm,J�k��E��>��jSP!V}���������u�`���K���{;�]������-�W�Ȥ2��ـr$�ľl�
0��E���ڮ?���������l�Q2y?��U����Wl{��Ua(�U������a�svqI�!e=�,�+�(F{��d�c�s�ѽ|A{���u������
��blb=O(�(�s�<��!�!�'к���\�� !:`�$]Q<�V#M"��Q�E��?	+v�����n�`]0�;(&n�lv������kq�X��ݛ��n�27���e��\O��=h*r��&Į�t�ˈiX���˧c�G��!�4I�!�HS������Ȧ�uwR�FW����ơ���n��3���h�11�k��4�,@��w��=�m_��S;x�c>��4zY�́i�K��űL�($^��G���	�y��4�	]��nk�~��R�� g�ʿ� ��j� I@�Bb"�:�����mrL�| �=�����I��'�O�늶��S�5կe�	���ĝ�)���@�#ժ��G�0�TR���G��� �p{��4��j�	E�z���ɻ���d.M���pXxٱ�*}�)2,rh�3	]�3�L`���\�� ���m!��#����y|�)��0%����"�3�O?��5��͆�
.���W0%cwL�i|i��HkZJ�4 �G��G�1�w�(\]�U�6���t��E���
�%蝬ZU����7�����ﶗS�%�b�����;��4�i�R�j�D��И��u�io�l�n��1�vQ�:�)e��C[!' �n݁'[z,�.����)�V8xu���\�b	���&��V�:�.��,���{e�*4a��t<T��}PTĿnqk����D|�1���*q��NDõأ�1ڇ6�#�cj���ȏ��
r,EQO��X�+���
\!Qi����|W��=�g,�q�CHF������2Zچ��Y/Պ��|>y}$w�bM�6821����`J��.}(�}���~�_�'z��y�?EfHI�Qv+M�{l����
��"�$XK��Βi"/sWc$|
�����^ב����\8�
Z!/��N��Dm�dSi��vK	�^b(߬`T��]#8鼚���Sx�Y�׬,U���1}>NLt�/�I�����ڰ��k�SW���B���F��^$(�e%�S���ɲ-
C�L'�E,�F ��o��b�����j��ӸN��
�o`��R�v� xe/`�5MQ�<;��q��((��i���㘀!Ԋ�D#��E.����6��+�����F+ּ?�����Q��hzU��t��;��w¼}GϞ<����a�)��^]Ax��͠���-��,����c�����w�QM��UݠV�/f�l6�U!~8XlxV16EB    fa00     f20�!���{��M��hu��;�=u��?�B��J&`E�<��bx�d]`��Ry�WB �ژ��% Q�wM>!y�滲�}�2-g����;4�ɟ�Z��v��Hv3��c�	��3�@�$��xm@T����C�d�i�L	��-�O�&��C�����X���Ϳ-�V�`^i׬ʁ�\:ph�9�"$s?���<mu���W�w?n� SM,SދU�e���y
�ʃ`�s�VpJ�W^%�q�i�3�����88a@Z��>VF-�{�O�bC{/�uP����"s��
l�E$�o�^�p��P��'�s!��ɒ���͝��X��G�Jg=6�0�Od�N�D5�D�B��9S5k���J�+,����DB���G�����IY��!Ζ���Y�M̺�s9m�Q���p:E؄V���B��`?���&rU�1�
-\ia�9��|���W�`:3����}���S�ڵ��wi�� �s��+��W��zB�г晓m�:����R#�p����U$��9�?�����)�,~����j���� �4n��(z��I��D��<@�k;���,}�P�B90�&�b��>��!+��u��˩C�d��y+#~��^�i[���ǃ�T��z�¹���.��4:#}���w�`��g��*�
{Z��o-z��A284�CH����6��'^�p]��J��YO��;�h���yK��N\3_�Y��8����ʯ��j.����9j�ȬJ�7+:3���u:
#��#�܏)���C`���C���7�S�l�aKYǒRq)=e�T4��CiߞˠV�c����<u���q���5���@���(��vJ	��8':b��h>��6P��O�ۉ�,�Ƌ�����8TL��>�/�_���x�5��r�R�+H�F�2����g��!J!䨲z����g��È�ĉ��"�{A�A�� _�h�_�k�5D��@��9�S*�fa6�7�)K3JQM�O�hk�BB�u�����[�v$��S	ƿ���x�q	����h%)l�9ն��>_����Q+Ywz�k��9Xz��-ϫ|��~����14o�=����}@�!����3��;�������P�}�>��`ϻ�P:if�H��&D�-����;~9�ş��Z��K*o[�]����N/!���'��S+Ew��c�;�^����)��^R�1��B����Ď�7��rI!����qN2��.[)�8;�n�2x���cQXK˝�z�(E�-f�b���X�y�~���TdQ�H�3�:�)I8.+��Ó{��Sw_{s�T5�ޞEn ��5O�c@�+���a�6�J��y����@$�m<���k���ϸ	�x&驄�U<��+3z���e?˓��I����ZH�=@�����(�0Ulւ6/����J����q.�H�����k�������OPV���Q�Y�9�vzW%w�4�HX�9-\�|]O6�4�ڢ���)6�r0B]��H������'\�άkǽI~}G�|'Ɨ`��x�S�ϯ"�;0o�NJv��I���!���"���t��o�ʅV��G�c����^�09Ө�\��΂�t���ïW3��ׇe���f�C�Hؼ�<�ȗ~���!������0��o�~�P�Y��;��3����Ka�ҷ̿5��]�/G�[_g�ha���I���46�s�wXf�H���<�K��ǒl1�x� �n����G�Ve+�8�	��O
�� �:��-���塓�7:���lTCL!��~~|Ss��5��wo>6���7+��/ha2��Ne��[N���K�}���&6�|XS���mfsh/�sy�c���%�H9ܸe=�a)�m����i]��d��V������V�Ph0`����<NFԒ,��+�W���u�_.(���(����g���Ԍ�l���֟c����h��o~�)m;�%��޹A���QX;Io"��!�\��~xS����;&�~ʟ�%1E#�İ5x�$9Ae��W�&Ò
� Rn��&�|�b�(��w ��f�՘H�L��ԳzV'�BF�&#�g���YE��~�u�����a��z��M���!�IN�M�?h��A�U�vJQ]� �uC���v�ͳN��AX�u<�\J�v��ԓ���� ���"Uu�����'�=ߺ��ziXw�D�\s!I�L(��MɇbU��ӂs�� �x�ފ���ڣ��Df$��4`�ځ�tڣi���K�\[#E�#�RB�H���G+��ez,�� ��jR�51V���V���޲���m#Jh�m�����/�*D#G�nE,��"�N��X%�(��ډ~j��e7:��x�u2	��3i���tr=a����0��=�J�Y_;��oj�Q)6�M��R��-��Ej�Owi:���W���ѐ2c�x�����t���?P~����y64���kTS�W��� U#)��������-����ŏ�P�z�x�F�aZdW�����"X�SqG���b/��9��*�M ��2��Aq5�smĘ{'C��"|t����ҷ͝b�z�����s��?��㶎+�&6��u��?���6���G���&��=Τq��4�/ӎG���F�KN�Em�F=�j��o��2bh@���1��.��S&~��fX���d��q�k����З�PxS�Y,�ƞ��B]G3g�l�)�:5&��r��<*�n�m��}W槃W�Js��ĺ7QD��!r�5�H��'�`�+��L��a�"PU\�"E�gA�O�ӊ���U;Ő+� �{O���-�����w(��΍B]F0�G��׍S�?��J�Veظ9�X�u��@�'���^
�5z#�s��>��NZ3F%����8=�����T�������A�����΁b���1�P>H�j��w���uG�w���A��:��u���EG�*˗�� ��������S/@8�p�(AP
�E#}��
w,lՕ,Y�?9g���y#�6���70X��^ �4KĠ����]1��Q��fC
5��@��Q���MV)>	����M|�M���Y;/�>ս� p�˪t�Z�.}I�����7�DYt��3��yr��#����#�Љ��o�h�C�t� z� �;P>c[}/��P���,��^:I�K�}���X��O/��ڗt��*җ ?5&%v]�:Ql)1q yr�|lt�ə�nAJ���a9��f3/��<��ʱ�]-e��la��%��_�L� x�ſ�R,���P6+}�8#ad��3��X�2w!��`J!ܛ�ﭟlY���� $�te�H�RS|�I�V�42۫Ĉ��zmr��3�@�&5�
J�Y-]�-d�=������欨�|+$iI~�ȫ?����1"9AA:+?ѝ���"�����;ҟ+�d�#!����=G�j_�B�Г�\��a�l�y+�Zjۗ�e�v{c,(�UճӐ�9�/�/�F��nIk� s���g��-�< ?��X�C��]�d����L�kHU��9HZp��P�*�ʯ�Q��q�bcP�J#v����
+Kz�|}�"�n����k���>�R`h�oH���Un �+R!k�j��:��PI�b~��x�x�ȧ�N)p�1��oq�w�ɩ*���O�/x��<�\L"�Q`�_��rc�� �D9�6?��@*g��Z�� W�K���pdF�X��g�-O����ٱ	�A`d�D7��W�L�g�r�H���w�-e�������-��i�BٗD�����>�����rh"��瓳���XlxV16EB    fa00    19c0���WR�^;o�B8�h,�0�����2�iGKH>)Ӂ(�bj}M��(-=��OTq��=���,rYBTb�Vץ2%~0k�j� E{񕥌*�j�o+�An\�]4����\�t&��h]�ֿ��h=$s�=̩�8K0ū=[�z��r���6�&Dz����E4�R�	v��}�m�i��>��> ��wM�vg�{���g٤��`�<X"��r"���!˰Vӊ�(���[0�Z�(���>�Ə�o4N�I��a&8b��h"�C��j/�Z&Q�&N~�r�Pk�/!�J����c�r�MC����į78p+��-�D��?���d�� ���h�ZS�2���v��)5��l��B��̈́�����s�R�rI���i��1D��X;�j}A�Omk$�52v� �0(F-5?�SV��޾�@�B��K��7�P4\�z�T`�P�)$-�ֻ��u��Z{�'X�e�]2���#�j׎�=m6xA���TC�:x`�:pE'��Y@=_�PQ�P���摹�Ja:�Cj���I��2=U˜��d������7NW�{����vEG���
�2�0'�\PpÎ��k\DkOm�t�N�"Ņ�.{�v*k8�S�-AÕ����{�aJ.�h��
~#�����PK�➁����G_�W:(�oszа�^"�H��/L��lo���o
hz��V���a�Η�_��e��ߥ����J�u�rFմ�]Z�T�m?�'o�ZI,����2O��Ǩl��� �3duO��L$x)�Xo��=4�V/�`|�9��_�*l9���e`���g�uQԩ ʠswM��`j�1���d��+;�O�kv�Ȯ��׊��ӧ{g��ùr��̬4m+�@����a�¬�}�V^�/s�,ҸHT��w,a7��/���iU
�p~�����E�S��_,N6���N��(���Z�������(E����}E1�[�n�f�5)��C~� Oe�8��A��L8u�`?�y�@�!Z��8��|8�%����I#��6��P~ )n�&Dz'�!�f�&2���(yV��q=��ྡྷ��O�G1��d
J2<<������t[KՑ��jv�0�� �_¬�/����[PH�w�ю��Gӝ�-Lt��{��c�.Gh|�k�42 p��n�g���Hz���y#�u�TǢ�y�{�؜=t� ��2(@����W�eȖV*�쬠��*"x,�^�S�ɖ�?ɹ���HԢ��6"Y� 	��=�z0���v��n���H�ý� �1��uQ��C ��^\[�r�Xn����/�LE=�I�SP�9���4i|T-��0��;�0���iX�����*���Ҹ�͸�QA̽��Y�[�G���xf�r��[����U?^�ai��6��V�|7����)�.�砢�e[���*z��`�/ϑ�K-:N�`ʮfd��ܨ)�	���߄ѫ�$�x�k����kE@Sj���9#*��7�^"|�h��۶e��_'yo��BT2��a'�TG�-s���֝�1���� ~�ߛ�Z�ҡ<�*��ب.���je���n�T��x����	�+��볦���\CV�0�P�ڻ�C�[�[d�)I��xSJng����p�}��zn$�`f��x�pŅ
�2?���)�;��G��_���I�R�Yn��H'��Ч�Wf~� �j ��ܬ�>5.8FpՌ;�@�\�^���tD�s���6�X���1���AZ�'�D,��_�Qe;�y*An20�+��&� �\V�j�0�pv���&z�"G�_dǚg7�)F�'��_� ���;�L����z���=��@$��)|��i��`��-|��uQ��$�E�m�>:� P�
z�̝Юt�g���t_n�Vbce�z���uY�yewt���s&W��)� o��+�r��pYZ�Z�X��،?Zzu�7k�F�>�]4�'��!2�SB�b�*���IzP�\��t�^�L1��5#d�oPi/7V��Z��ؿ ���z��\���B�ڑM�Ɍ�c���p4���9��O��<� "^�'�N���ԫo� �/�/c\�F�3�1pR�W���ڼ���y�t�3��������F��E��d1�6�ӆ}B�Q0�+%\���fpf�P8:V����ټ#�GCi;̍ai6�U���u��	��ܖ�|@��u�9j�p�1�P��i�:T�_��;L���|1_��_a���Óɓ��P�W#Y�:�T��An8�����3	���uC �Oső7$&U���#shf8P$~�Zo$� ��AF�À:�=h�d��d��z�T����n�iuv��|\�����q��BA!����q��=��l~���wk3���x)�Ubz2�e�Y�a�٭{T�"�w72w
�
���
��GD|�ץ��  ��70)�nW��Jx#P�B�M�%�D�Ѓ�`q���ID�($�E��Xp�<Pj�7\J�)R._F�q�2�7!�U�ݍ9EyE�&�3�rio&���xR.^�s��8�PQ�u�5�Pb��ڬ
3�ɜ��گ�n���?�Uz�� O9�i��������K�������\.�A�,���jD�>� �˰��cI����]㒈�c�%߽ORV2W������ȩ�ٸ���ȝǖ��_[a�S�vd���G�=ף6������&��d�n���[g?��qA�i��nWF؝�>��2F�V��^��<�����7h�Jz�A!���h�
�ЏT����FmF�J}��&muW.���H����`b
LCH���;����6��z�;�<rx���Q>4�(bc!�����>� ���n�W��HO�)!��0;zE �:����T|�����N��h`l�]�����hK��tϡ�����N�Ƥ�N��>��9d���eB
ݸ7�V�+��c�DX
s[���`]`�Q��FQ��k�y5:
F2-0�:y:>E���\~�Yמ)ڞ����e�}{8Gu$euY*aa��Un���V���~ތ~%Gick�U��Y����6*�+M�i�\�i*[y����'�GU1�pS6޾V��~�E .;V^��b���}C^�7N�%eG#����_u&z	4��ldx���s�ی�,|W�ag����>��Ў��E���|��Q̺� ���������gX�I���y�N�/����`��QCz�,}�)��u��{qp�@��,1]�'�+�~�l��2N��)K5�%Z~�od�K��a9l~YH��4չ]۸���Y�
-�_E`����ω��,�ԣ�#S���?vu��e��º
���o��P�LD�_��:.��h��Д��W7�f�Ψ%��+�K����St'H?6�<�����w��u�Z��
.��fx��MSoE4t����&�T���Ţ�*��3�
�A���"���f��4�E+vS����R�ӹyӡK�8��_k��B�
ם[�5J�lT�ۖqHT˓0� �!ل|�E����Gs���9rC΃G������R����� '5���U�.�^V/QKT�5Ճ���_�n�\�%���(O���qysؤ��j^8���2�0�:hh3���Y�BT5shQ�釔QO1���̘(p�[�>��<�-�}�ݾ��s���Ɂ�=�7��&�&��b���,Fj���4t��l0!B2���{���t� z�yx��jM/����|��}��EG�w�z$z~6ȧ^q��R6F�tZ#��G��!���8��A�ckc�dI ����S-J�F��DǢo5*8H!�|�ո��k�m�9o�nЭ��Ć���� ~�H �rs�?��n��l{���pD�>����'�S��.��b�5��d�s:Lf�XhD|�)� l�h���:w��� ��y��9G�b��F�Sk_N#�xW�A�Nɘ���T�'��QOUk��t~���䌿O��~�l��!�%���R��t��Ed:�e�>/����V���d�[㓸��O���G2��n�FyS�:=r�bk{00�,�Ȕ��f��D�mQ@~����)�M\u�B���R���
Y��hl�!�k��֦98>�� ���`�G����n�U��_���]@x���	BT)7#��;x�.^�lM&]I�uIX3i��;�O�z��V��>vr}��t#�.��l9ͥ���'a%$�L�]6�ϭ2!�̄���N���¯[ސB��3Ԁd
��e�oc�GFt��U�j�2�}'�F6�%�'[X2
` �3��L�r^��$�3)�ӎ��zVVEm�H�'�%���>��K_.�}��@��/����g+f�s��,=������:�e�ʳT!?ϻyV	秚��6 hC��a��L�Mo�8�1�k�@*�
ӗ�+r>ZX�8�}Z/��W`_��^$wl�u��-�S$��(��a��{�w���c�]�Y2%tB#ِ�"+N��$s��,�֯�:��i�����f�W��O
NS߹)�( g�L��Q�.���|�/f����::���|���,�Gs
}�	l%��9�T3,jU����VL^�ߖ�h����i��]�Ztt8�ߕӉ	N����T��� ��gH0�=W.
Ã�-6$Fy��v�x��0Τ ź�����֖A�療�o��	7謁L�$x��-m��{����K�M ��F��c�t4�g�>4T�{�4|�GJ{�s�WI3`F��q�l[kvd��A��ÿ¥��Q��{�-�6n��b(���ջ�^� ���A��<ufV]P�e�V�ꍪ���k�`�D���Gc;N��#������^��ꉡ���LY�I��4)�J$nKf���?T���k�:C-�,hx)X�\��+����A�@�0�>�L�mJ�hKd%2�
��:�4wwo�
�!+�"QVO�3Z����������z��u۴�d�3M;6c����wi=g���p�-C�d6�<�D�6h��kA��uM�*<[�j��VN�oG�"�g{ K��C5��� ��D�(�F� 6ebO�?J5�0�ny5o������jޞ-b�S� ���\��䬩}?(��l�|- D��F
�,��⶯R�یmw���"<��fS�+P����Lv	wIzU��눉y��l�!'�'��+O��&Ƥ�4�kȦ@G[�;7uR��m�,�y.��?�G��XD�#�5cz��*f(���"�	W��C�p��7������į>ۢ�ţd���cH�b\�|h�N	�@q�?�z��No[��~ �*�����V+N~��]�R�'~𙆷����@�)�M��;(�:/��*;�*Ӭ���K��Nv/�;Yɾop>c��G�)QV3SZ� 	����q��*��#KوrN(2n�Z1�_��Tb\��
�y�$������V�֘�J1E`x8aS0-V/S 8 =Kv����â�g�c�>��A_-`C��h��v�eB�-������mke�NJQ��CL7 5Բ��s� �ZJH[��P3H��'�CF!q>���3��o�16A��VC����y3��P�I7��-�p�����	���$˄jO!� i�Z���Z7�<.��#C��na4fh�R�z~	�0u�N>DQ��=$��E
���B3�D%�5T����r�Q���b�[���sD�V�M�����幂S͕�.<E/��=���UfM�]i#�D½����b�ͩ;�I��������@V	,(�o�e��.�]>o�Ȃ��ZԠkoJ	�-����z�Ǭ9�Cc�� (�Ƴ6�9�@J��m��뎊�.Nȵ��^���9%�1�������F�.Tl����u��,��S�e�����-�1A�N:˱�@�a��J�IG�kA)��J;�S�3s�]�$��e'w!<�<�<����x�]��)<�}��42_Q������Zl��Yr�261)�}A�!;��G�ք�Q_8�0I9�
��PXt=ڼH�ӌ\]|�_'U��8&t��w�{���u'|1#����}L��êm�E2�=�&�`I�-�l��uV{?���
�/�?Ð�~P�`�(�-!��uN��I�4��rfL7s����S�������	/Kx.�h�WlǴ`m荕M��7�as���+�	����Am��g&�������:����аx]��G
2N�F��-��ڏI�z����tvJ`\d\R��0�I�x�|���v����L8��$�������<��ėK
���p���:���`��̉�Ӷg������Y�Hb����0���ck��XCv��U��^�v5�y?���hD�P*n
�ה��y�yA��q��*�9����5�\�.i��������"�/q�"]���Į{��`FD�/a
*��Ml"��':��7q�rE7�m�r!�[�m�Y���y�%p?A`�᧢�NFXlxV16EB    fa00    1ab0p���Y6s&�~\Ұ�~�nt|��2�-����M���G�������k�mO���Y��a��,�SV�m s�X�5�#��L������Uw�� <{�Lc�:�Cv(��D�%h�K�	j�>�Y->�>�kO�c��{�] ��ټ�Y��X+�"��ɐ0ק�%�"�q71ع#$����t��4���D
"5�2Z�^��hwf;����m)���Ps�����q����{��&\� /&�Ө��TM�"k����/S�w�h-��;�fu�&w��Z덹.P^���5���XS\� j�i)rV��ʄ8M��;����7���J�_�ns �U��Z"P�^�.��ୣ�N�0�L����1�*a^4�<0�3����f�����f��y���ȅ��'DW�=��>A��Q�}zL0��r�T;�H�d�%��h�s/�Sg���Luo��n��%��*�{�n�U�$�0`�~�/������z��2|m�c���P�����9�u�A[����A�����,�j-�-��vg��?l��Mv����wV!h����1���i�g���G�2�+�e���\��~�^2N
 �,��R<T����yρ"C������}Dk��b�Z�.���g�.O�e[;wή�Z��E��m�o���f��?���}N�isb�r/���<b��``�7
��4���r����7�R(��}�o�_�����wS��mmM�'�h(d��=��(�L(ox?�3�f��M��:���I��E�fe�ʙ.�Jx�g����-��b4[�)�Hps(��av��]Y[n�U[���x_U��{M�jK֛�e��皼���<k4ʽ{�� OY �qoj�W���l&�R����;�9�#��2�~�j�c3F�ǝu������J8�K}�h�a����TJ�-��G�aAkvL� �8K@���'�O</��[�L����;ȕ�C��B(��	��w�^~�t�)�ՕW�B�&�[���
�<0�:�U��Oie���|m+���~�=��[O��FV\����Ʊ�s������B������tm{�_s�M|i�99����dZF���gSrb�LSmn��N�z�[�p�[���^pN߁��W�'������3\��r���.�e`�=�YLl�]#]C���G&KA=��wD�p=aÖ#�ȣ홛}�����x�"�*�~�9�0T������i���f�N�x�dvQ��
���t��z�@e�$[Tl��H�m�]n-H߹���xEYGSڇ��~|8���Y�K�i�-�!3J�3)��]
�2T��P��
H�p��;����Ĥ��f�7V]˚�P���-	�W���z�b���vQ�<rʱJ�E���z���[����Cbw��?������)Ӓ�,!��G��ϥw9t_I���Á��h��ĳ�.�rWrb�m�4S�XO;ŕ���M�.��.W��Y�:R���!�E��Φ�#����E_��yC�����1�E<k���1���k��I���tLB�Jc��iw��H���пh�㘱�E˔�1�� P�YEN��Q/��Z�	����e�]�ήf���c�rp��K#�Uk.w$4p��N�T �+��@,��7Bۿ���@���uѕ'�+��\�\P�ɼ[+9ףEW�ޭ��e�i��-KS+���3���\&�@�ͨ8�.��E��a* G/6S��Y���O�,o���~���EM�ݙ� G5t=#t����xf	�4���"�wG��4/�kb�uZLf��� ��"B�R�p�)T�����pp�[8]B[䗶�t��x��Cw�MC���f�	v	��͑�Ȑ�C��V��ɴ�Nݦ듴����ͺ�T�S��՟��k��P`�R�R�~��>S�K�bIR���0�j���\C����$�����!���t1&�`|��7NRz�k������Tl&�r�Q��J����5φ@1j#��Iڑ�do�%^��;)�aϵ�e���9���1LqP@*ą��G��xr���lj���i��U�sڙ��4,��->?y2y�T��X7e��P��k?�F�j��t0���"hin��F���3�c��;�rm*)�4E���i6ٴ9�-f�{:u�ڭ���	(#J���#�ڇ��GlE���*�������J�ꅉ��/���������=���h4��
�ʧɿk����\��sĸUx�Q��NbF/X���c�`�Jfر����':��͛�ڑկd����'��C�5��	ŉTJ�J>j8��ؒ��2�C�Kc�*.?i�։��P�m7"�@bEP+�_ׇh��A��#�G0�#�,��o����̿��B����b�C9;;M��"#sj��q������Zk�`g=��I���E����Nn�"�"���4
1��SdWv{頼���^��1~����~ ��	�	�?�υ�X6�f��z��ծ��?�%�|9~SX�n2��\��� o��g�Z�~��$EkVz.cdu��!���}�� �8�ZǓH��KC���ٱ��\J��{��������c$����3�����9���jhj�ړ��lM���f�&-n$�GUL��rM�ҿS��� �}R�f�ݩ�^q�ọq�2�O/���W�����g���C|�?��	�
�i�)O�Vަ�U9�l��+�N���F9!��2��#��J3lC�0Ya�B�/4H�"j� bi�Ml6ӕ_4��	���B��Y�Y�L�!��0�B�߳�2�jтjߑsZ$hàY��[�W��X�D���x�{Y5����1I�^������p�����U�v�U�S��S�X�<�=��5 �������r8�W�]�rF�q=M��Gb?���gუ��9e}Ԉ\3#)4�w�QF�Y�z����o�*'�;�I��׉4��0=9�cCq���v,{�i*�숃q/�6Z.�|W���Ջ�����W��U�:x�;�#i[QuܠP��O[�,?V�(���@���u��#��jz>�r�v Ϣ��TI�zMh~+��'��˰V��ᆤ	�݈�w��c�cb�A�0i�E^���9� 猖d�tÖ�I�i��W�axL��� u�jŬ�����I���F���Ͽ��ņ
g<�r��것��t��7|� )�XBb�PWq��g���U�w�K�1%[���E>1>$Ѝ��e����b=�ޣV�v5�Ò�Db�J-�z�?B�K��W�Kg[�: ="2���KS	���U�4�Q�N�M��h���]�����a�7v��L�Y�9��}:G�3��Z�A���|�Cr��"��(�&�v+����^�T�1��*�x��~���F\'R�\�-xU��
=ӳ�T�r��'�F�@|��b9���PbTiX�v_�V����_��tQ�:p��zmS�w&�L��1�:ƞ��ϣ-�� N�)M�~'֕2��fQC�����jz@��K��)��B�>�t�ƴ�&�Q�^�~]d�Tة�b����?�=�/	
�X��M�	2�6Mx�QF� s��D��\C�Z��[�=	�ٟSzo�>_M�a���� �R�3����7���T>(���2�� ��vA��M\��� �s�j����65��F�:�����ž�B��"^�b7B�G4^rE���]�=ca����p�`��\���6x |#�������-�k��W���i��J����w	��.�4�lp�D·׆.X�nL�9�NC(���`՘_�@_|$��?g����M�k=��?H�;g�����4���޶)��ܷ`�G���}/�H�0�������(|h� >U�u[��",�>�AS������&ю���N�=e�%���+�m��5�y�
5:��8����N&�vҬr� ���7}|�����j��f���hj��5����M�8x�C���H�d�KX���Pf��K�r��ru���i*K/&��I[�
�A)-��T,���,�����σ���5w,v�B��Qs�%L1Y�b�'�S���%o�_�	g�T�cHY�
�Մ�/��Bѓ䙿x�a�X�$\jɉqC��t$a���L +,O�ݟg�;UG3����4s۬*{�Ex=����l���wo����
n���{�2�̷�,.}0���a&��;'�2���n&�v�R�����f#v������l�.�'X�Oۀ��Ῥq�J��cS����>���Ɠ5�9�U4�5�m �#�V��&3�l�ǔ��H^��y�"����O8�W�`Ќ�6n��Iȭ�ꅟ43�g�?�b��Ӓ��/�+0g�4�; ��(�b�F�B���x1� M�ut,�*�/gHxL�r��xYb�sL3!E��g��KUeM��&�������m��?0�\W}�����6iS����sa!�Q�H�C0F6JtvXك'�����em-[��-�/��`�Tim	@��p�W�L�1�&Ћ��a�1�a�ˢI���$
s�멀�n(��P~�ƍ�l�a���р�g�fLns4�bWJ���Մ��pPv��O���wX�vlkQi z �9~D΢�E�:\��4Ī&y&�ɦ��G�OᎮ9�<˱�l��\B������ˁ��$�͵iY�� :�ѻ׀"gC��y��pCv;�	�Xe�
���2%q!pSe��y��qy ���Y��[��B��C�	�� ���p��_{�9ܹ3=$�����W���sP��������o��9�32h^0?�+�)����X�\qJF�eT�ty��	-�(���=fWѣ�Li?أ�������$;�ϓ�)�qy������_b��w*�����"�(f�I5y�I�KY�@Wo�:�w�_Z���"�$�3t\���	��f1����$�V�$U�d�k��"Kξ��9f�2֏%L�Q_d()4 �n���ƽ�&:9ˮ��A�siER����#�MmUex���BUd�����'��z>)���H_��U~#��/h��rSrT mPք�vt|*�/����s�з�EX��O: _y�2��?���#ֳѪ�W��HyU0�#Ȇ~1n��F��_�}.�3�E�`l�����(Êy4�HK��>Q��gqa��(H��H�!��@�^"����0*U�~C���pJ�K�����v�O��?���u�0N��KCm�kub�l�� hx�z;~�ּc���1�'v*�^��.��=�߶�Z)N��M(/Qm���yhT菀��������)���N�R�7 ���U�.l���V#�d��Q�3"�py,�zθVIF���?�ފ3w��4�ݾ�5O�ԡ�u��,�P��Y��m&���m�����������ʮ��,�w���oYq�Z���I/ϑ��r�۫W���x�,�Y7I`�`@��=�]Tk
�Ș5�plDJ6�'K�N�Vن$"2_8j�%f����Ra�y.��E(�?�R��5
�yҭ�V��"�g�����l���R2)(��6#WJhb|��C%����pKR���[�K�n!���HC,��3J^Ї�s�̓��= ��jy�SI9$����^�V�xo��U�gQ�#����0�7;�ԫa��`YVe��"I�ܙ/h���P��_7��7���*�9��Y G䄲Ў�U�z䮻�����6�i�ځ�,��T~8�Zt*J�dnL%m�B�
���'���82��.J�":-�29�2�o)d��SXv`
.5���*�"5񲁱,2�L+���q�{0d-b=�>��壍�����6�hfxٷT럦8�6����0P�S�	� 1��n�|�N�V�0?d��ر/���K��?z��
�2o�g�7����
��.!U=c"��K�i�E�������xjr+ˌ(/�迉24NL��Q��|-f_�oq�ݔ�՘'��d8
�*tEr�]�7?��g%��-�JV�{�H�$�O�7����8֞1'�lx�o%zƠ/�C
P�_��>yA�h.��b����v4����n$��w�}tɲ7(��8��Aa����7Z���K�-�l��r���h����@�U]�a0��WZ**T[�?�t|������'o���i����Eb�>���mya��G�1�!8[[3_�R�����tHA�a���z�jM�:��7� ��}\�Z��d~�uͫ�|�/6�d�X{�e ���������eǙd���o9�ō�:Ζ3v��,��������J	H������ W�����-�R6IN	Fs�ВST��3��{�2��'�,N'�c"_g�n�V�F�X�F��C,ͷ����rd� O��ApȽ�[B����rr[����[=>_�+��\{�=� �'��'�<�w85z{m��\���,���N�imE��a��x��L���z	+2��y�4t^�P��b߃�%�do�Y�R���� �$�p�SZ�
�U��P�ޜ����2��}�MS�L<W�t�*W��*�`��G8�
��/$.�{���upE����gs�q|H�`�dh�"����2b̖U���"� )�18_6�(�g��fZ�P� �� *��L�ãO�{�#��X}���J=�`9I[���0T�A�N�W���>t����Z�ôZ��*!������I����&1��5l 'Qd��8e�1��D��F�a�X"�>;^�"x�*���&?D��e-����V��j�?D������|"\XlxV16EB    fa00    1ec0��w.F0U�y�̯PMZ�y��\������xH����~%R�Y)������	E�Zޙ�P��T;٠��75'�T�ί͚���D}�� K9TZ*�B���+L "䄃#YN(/v������]R:H��v��f��61$8��Ղ��$��$��U�o�S�r�e@A�Ȫ�l/�}z��ːGH_U�hO���rW؁�D�4e�#���)|?BV���2�m,=�߄L wd4 8f��!.�x��S'DgҕSe5�X3e����Q�3�������~Rr9[�K�5�Hw���r�]�9�u�`DW�]��p.b��`�)�x�W�q�q9�S�}�83(���s����Ѽ��\��ԸEt	6ck�0��^=��r#�W�M�?�ۜ��f(`��DQ��zŤ��+va�/�����M�CUs��=�ܿmgVwKd���XwA'�}º\ya�<^���+��3�N4�nB�{����?5E-��& 3��4��I.���l�W�L<�-w��'����LR�Zip�=���,<e}��7�s�*3xuQE�G�o<�������s�N]j�VUˢ�Y�t`>6TA��Uf�C�j��^���|.VMX�:#bw�"�M��j��^'Ď۷<���1m�	�3.�s0Drr���	Duc��~��05[q0U_I͆=)G)�o��n�ELݿ�~Q���k.σ���zn�v:՘Q�a҇�$�zQT��8����wl���4�k��	%����Fr!H����%�q1����i3�W/�l+��}�*؊{Q�����vL�!�`B1�_J]��רFE�����/0v��k�3����0��l@o��h~��S�@!�7᧢����:6���h��I?���!t�G�8�z�xQ���m�ۉP��%	�^�<��(��׷���Ȏ��,;��?N;2�=��k�/�t��7?N��L�\���E��Kj��*G)������"��@��-=��4�M��P���XP�FUߔ*�]���
�E�3�� �.(�ȷ��x͹�F�o���M�C$����P�9��v
f/�3|���?X��x���%�&�{���w�nB�\(��J�j2����oӝI��_�Z/Jq�mDc5��d��'��pڀ��\�X$������J����TLq�$�a���� |�S"����f.��q�b�����a*!1Ɓ}�B�R��<B�g���f&���|j�l����^��kJ�m2�׍��h���a*��jC2�)0H����L-��Qd���'4��yo�<�U�v�S������I(�bMI?e����"��ȹ�Г�I�f�#Rj�R�{V��H�U5D�Ul�ڋ�xt�9ss q�A/�5a���m���C�g߬Ia�m���2��t�_���&ʪ��M�ē�oT���{t���K�z�mMȰ��W��9��CP�/6���X����B�Zr�誱��1Fc.��2XP&b͓��
Y=�O]�p���u��F��R�=:�M�~����9��������� tKR��\^)qH�j�rw�g�r�Gx�t�>|�?|+���Y�����DC��_KE���.(.���� ����S!È��W�	��T�N���@D隗��yT6���I[����U՝�S��l���C1�௻l$1#��b�}�?�G��,J��
9�t�~;�}�h��o<&�x�Yk!�XH<�	��va4_�ߊڑ��ĉ�7��ɼ���[e�a������� ���;�P�?�h��=��r�Ëh �Z���}������vS8VQ5VgO�^����\A�rh)�	tG��TM�
&#չ{&�}�yd۲s�ߔ�h%����C��sfQ\qga�+�s�T��ƺ~��i�kN���(�i�ޠpA>��ݾ�<g��
�cp:��|����� ���L��e�� �`9�_�CN�\[1�[0@���u�~91��?��@,�0P�X�$RB0+жkM�Ul�C\�n�f�ğLܪ~V�~�5���;!״�C�9���FV���#�)x.�.���4�1�����X<�!b|UW7UJ�9�9�{�5�P�%@sBīF~��G��$�0P�ztw`����'��
�_0�r�H������]ɶ"!� ���Ù�0�[zW�s`7�v�-��p�J���7x�RZ�ۉz}"A[>c�iT���m�p��+{YYw����:��XSA�Cp���J������tj,�4
�j�<�{~c>�sRI�%j"���m��sn����4���X��RШ����}~Ab璨M�W��N��<����n��B����^��ؖ���G+l�����Kȫ�=��_mp�u=���vi)n\�7�����B���9��gC?;�́_�f��d� ���x�^�;E�!2<���倡��2��q+�Ϯ���\����$�АQ>9�A���2͐6Y����a��7��`���9�*�hK��4X�J=_��5��r�^�ڻ�iw5_�D��l�K]q���VT��r%�8Mi����="�x� �@��|Op�T��J���GZ~���k}�3�nj�,iD��9R���3����Y�^���"��ט�Q��J�O��Ę� 8g�W�HF�SiQ��G�h��f��� ө���buÓ�7�%�6'�S��w������?��}b�^d�{�	����v�l�lKԁ9D\�ܟ�9ͫ����ԃ2(��v�,���~:4aA�ݛ���}�������ȝ2�h��2XuڎɈ]9f���_�@��*��⟡`��7ex|+A�7�G�RE���oȴ���b��KYfʭ�X{1��B-|�%s�?�̧l��;
q���5<�X��ݍ�j����$�+"
�G[���m$V|Xx��~��T
)CF�y�N��$��m��)Պ�|!�R_����YL �����C��*N�����j�eQ�.(�bK�ўGgeqH�J>^Ѝ]�� 0�A���0A�4�Ci��iwK�p���Y��^�$�%�r�F��6ڏ һ�?ܔeaN�U Xr*���	��1�1��P��3�C��l����� 9%0�}Q{d���0����I: �c��2t���\~S��iZ-�a�m|��T�����^K7-_��}�\�Зgi�e�:-�Gy���/ZgI����,��J���;8��4~���~���
��V����j(ʯ�������ӏ�l��h��4N�P�o1�5���߾��Ȉ�ć�&��~+V� �s�Aǡ'�0=}�vK5R^Ud��N�w�{�H<��}��o�
�ؓc�7:�C��d,��\�8���ì:�����n�?��Kl&�+��s8�i��`1�%	�aN^��uç	�Ӆ�3�A�Ph�wع��1=	��I�K1�۪�� ���3���i�ށ�x0��4*����J�5i9�/\��"�<�]4?���s'zj�o;�s�5��*xX9��qbYNoU#c�Q�2Y �e;��A��rj3s]>��'�>�+&>��.��N덋Ai^��<@�č�9�AW/�w�J�W�,�`}��ym���$E����=�
���C��t��[8�#I���Q��I�܄�c�_�J�_��C���λeS�l׫"�9x��y®�
��q��Q#6�)�ɽ B���Ӑ��en���s7�:gt�KB��2�H>��8�$�5�I_��KVHާ��	��r"wt8��|3��
�Q�6����qB��Oy6�ً�9��ȗʝ����Ǌb��,JKzI��m����kA�H�aF;�N���/t�s�H�IS��!��^Ä�[�W�S�h
vp����
@%D��e�B���*�'"b<�l'��G�tK���N��Ghd���v1Kn��Q?����#�ڹc��,(s���`k �����k�(����[n([�܄�T� Y����e4MN���и+��R�GX4V���a�c�naY'�S���_����S�q�_����E�����G��pulk~� �B���0"j[Yx���P����� '�}���%i&��^0E�I/�?3�)8W�␜!b����
�.L���#�p��1F��/C�mC��;�>��[��e��)7q�;|M�J+���/cJ�6a�&��	�� ۄ0�"��>z<�Lغ�K"^�V�}����{�0(�|`�D���/�UqCWA	�A�¾\ ���ݏ���2����y�o�`$����[0��*�	m��]+��l"5���5�w\P_It���V^ʤȬeBL��EG����҈(����ʨ�9��(g��tTdy3у/��H��m0wy_f��b�:C���u����=�ۯP�����fjҝ�y
3��EқA��˄��b�byO5�r�7�hQ�X��)�мX:�P�Z��F��]z�]��C��A���/��������������Q���w/�O�UD��DCܬ%�l��}o�h�۬1�]M����$�X���T��:[�Ǻ,#X;F�e/��{�4R�sϽZ��hvK͗ȑ��I�%���	��F���'޻D�T����v�gQ�[�k��0[C��=�ፈ#�Z�,�/\PY�q�{��b�>�ƙ2�*{�@�I[)Y��dOC��25]>����8����Y{���	=8�8q�E�W�A��F�+��j~~T��n��)�5��E��}j۱KG�PU��uB߼��2ttcC���6?.6&��V{�zWQ�	Έ3;oZ�׳Q�4��u�B��M�����8γ��o�F�����'J��-S�+�9�KءAA�M*_U�]O���gK���r���?[���l����〔j_l���kUP�t �!�H�a��vP��-������:���b�&#���R�N����Ko[B����{����KJ�r��#�*%�a� 'R A2kv'�M������q�B���dnL��B0Eߩ��9�>��!�6��O� .a��I9�@<֚�S7>;M�^w�t��~���n<MB�L�vPBc�M/�����ț�Hd�D�(_�C*���B�B�aD�N�P߰�H�tw�[*-���H���\�FMB�������: �s|ģ����*�D����7DU{%e�����?ch���O�ڎX�u����:��}�~�r�)�	
���WnI�t�»������r��I��k����07��Q3�i@�FC�4���6�j�[?�	�Cw�����V� �c�EGx�!�x�j7ܘa#V�X�T�&|���u�O)���Qg��~uRq��5����C�?ƣ
S���yE�?WU\i�w<�Aw�J�Dc�\���E������\����N�sƧ?�_�(u��ԫ rs.�|g�?�Hڣ�L�z[���;�^jʚ0oF\#�t��S� ͇��Oq���:�ξT��D�|zF���Is�s����"B�R�x\8�̉o�~�l�r'��V��̡������,�[�M�a�p���4�@"M�8�^�����W5���	�ʏ���]�C�$*98��ce�b]�)l��v@��Gt!z�^؁�.�/nD����:9��_������/�7�Z5mٴ��Q_�ȟ�̶�r�Z�U�f����Ņ~�s���&�`�wc��=�f��1hH,�h�	io�+���~��(����5�XFp]�T��;8����N��Dr���L�>�6����
w��E�kuJ-���1��0��z���p��>�AXU"�)�*V�w&?�;o�(>��w���R� 1�}x�1L�M�aby��AЖ?fR������A��P�i��kĞ6Dj��"�H�ͮ�s=�WW*�0��A��r�G�1�qU��A�3�`N\>C�+�ef ��W^��2B��ΰA��z�����ꮨ�ao4���1P\��c�#��e�qn*F;�)f]�[@�W���ʽ���i�A��L�d��A�LIG�նϤ�>jׁ.�/7,��M���i��iWh(C��%P�ɨ�Gn=�T�����<qa�H����aTEE)Ÿ�Q9T��ۭ�'��
%13$�_�nK�6�K.2 �XF$71ly���T�W�sˎz`��v�nO��m�S����)���z83�#���.թ�]�K�W8t �M@m���7��\V/�M�yQډo��9;<>Ld[����XC����SbLrUZ�1�3���{����5�n�:�e6e)��vf�������
H05�8�;�8)�6oe�LC�a=�'܈��҃}�#s���3��B�)R�᫲C���=��S�}_���������Ȥ�Boi~�I�K�׸~@�+�TmK���ۼF�_=r:p�Cخt"@?;c�غ���i�Z��
οD<��8�����S�o�0��.=�X�Uͧ��c'��>��&������W�ZL��~	Ni´%T����&�NxZ�v�9��	��@[V�X��d�(י|����8��W������o��S��ƞ�c'�ne1p�X���M{���=�A���I�:)�EI�Z(lk,�߰�h��uKN+~��<�@��|�@��^�W��~�._�����z���iw��K�*@�!�v�
 SL��_WN�n��6Y�H,��қ\�Þd�H�!�U�)�G�	�H����bq=Ԯ���S��|&��)����4�P`�vB@E�8p�$�2�KSl������sWd��K|��_���)HJw"�$��)*�*n$����x�bGW����d&�7���h@��ۇ5�ZU��_^/�Ɲ D2�Q/�=�i()m������I�[�P��"ܯʑÔh�F�ɛ���ڙ�O�'����,�IJC�QoC1Ҍ2<�ߔ?���,Cp�<!�+4P]ߒ����(�$�����HI��Rf�V�żBW
h��Bչ�����aU6�p_\	2 �vI�F��鴇>�B��DH��խ?�rG_����a+E�P$ӭ��:wYkp�TF�ئ��k���l&/������c����jiH�q�<�|T6��%*X�BW���-���z82�γd�CLU��-��xx��g�6��?䵠v��X�a��±�ʼ:s�Ȁ4����O����:���F��U$��Nr&���B�	ȵ��FP4kd�Q�lf}�FgUi�쀽�y�U�mQ���=5[��7D1���I_�L㸂�����1Q��]�˜LpʱQ�
�l �i9�P[SW����r%���GI�[�B��RH�U"��w�0�R�G� d��3`l�΢���N�D(����1ݩ0:��t���8����1W�-���ʰ�Y0��:;Aa�ͤ�K���!vPl�x����G���i�3�8D����߈M��t~�U��J:��f�K�)�Q��D����Ǎpder�Q�B�B�O���o��}�b��T�SE�3��A�6
��תz�Ut2]A
��2�&�n���ĽGM�u�ћ�c����7��8ܦ8!<����S��/��XD�f��Gb�t��,��kx<���SrU��'d(��ʪF����$���_'>2&6%��B��VS-���,8�4G��Յ��kS,�H� ��t��z#�B���՜l���p5���J��:ů�'�E����?AoU����.��D�b'[ޖSB����y}��Jv�:\Nr�t���.Ǉ�ᥢcJ���Y͠��¢t}�v��W�B&Z6����V<l���r�Q}E%�xs��۷�r^A�)`�����N�q��gU�*L�i�p|��H�B���nE�) 2�)�)��d�
nߧBafXlxV16EB    fa00    1ad0j?����/���r�o��]w"���q'Ǣ5�,'P�5(}P�X��}�DIcū8)ĮW`��K��m��>\��
���X���Wϝ39�>�W#'M�!@j"D��ܮ�g�y�V�#�W�L���Z��7�&�M��׾%/.�b���6�u��������Ԥ}%m�X;�v�)��tcV�nSU�]k#K��'�ny�*��_F �6�C	�2��5%t
pJw�����̮��+�a+ݶ�0K��x-�#HG����(�ȟ�Aa�ay����~"k�<��f�bK"i�?�{���T0}��������c��j��XE�9��5�"��:I�0�y-��\��H5i��{�B*��em�Пg�NL0�&<����n�����d^�| ���en�^A�]�I��!�ܽ8]e�Nz99�|�-�c�壦�+��u�,6�ͨ�k"[ ���E���Cv� �6�'��s��95P�B$0��g�lpx�J�z��s��y�.W�;�!�ɜ��|����}=����� (p�@�N�»����T����4^�cfe��d��(WKğF�u�-��NU���s3�l(�ݱ��*�n����2y��u��"�\{9g�-�RmC�<F��,*̥&-�d�}k	%{�N�9F/P��jh̬�"2�Nr{����5iЮN�l�,���J	�V��+�6�����"Q�6紮�'�X���Z��Tc�ݙ%)2��8PV���jR_IJ5x������k�3h��e>�doYH���쟜*��з��c/ၝ��2�
���ea��Ղl�PK�ӣ���� ��m꿰q��S�$�O����X���+,�����ԭ$):���	ˀ���M���|�[}1�<�S(�γ�'?P(��RVm�6��UY�'
sk��4�}�2�D�]��l�m�%*�쭤Z3�+�ƮG��>�C߮E_O	�)����_h���d3��k��C�I���M���u��qô�;������a3}�;��Z'����e����8�W1&$7�@���.㊹ߍ*wI��:�Y��L��H���M�4��`���0Ozos�p����+�
�"�_c*j����T͐<g����I�L�y��a�DvoE�F�������O8a�O�by��˄>r��8���+�c�r�<A�����K$����-��nG^����I~�b��y嘿�^Ϯ5�4k"Vnd����u�w�E2���x�O��@5�'J���0�0�d����s�� r�`H:5΁���� ]-t�t�����Y��/�/���}�t]PG�ߴ��m���B�I#��.R��h�4g6�VW}*^��܇�rT����Cq&_��2�O��ڕ1�?��BB��To�8�.ol.��x�m:*�c}����w!��O��q�`7���f j���wv�����6��}�g��S� 8Un8��<��'=n�Ӡ�C8�NJN�*_f��f.�H�S4/�g�)�G�ο���s���z�B�?�f�,�R#������&Nr�"�PU JG>�Bj�Q��)ӡ׭�q�=���z��aAi������Ji*��T���H�g�J�oYigJ��YV
�h�a��ѿ�$�렲\���aL���{E����7����=�}���X���y*�2�7�E|����r�68�p��{��,�������Z��*���(܇�2���9������?�̣�C`�QC�����A2#����B���#��nF���*��� P�����NG
~�',��>�]�F��R؁_��yO8�3����.w��c��t�A'�� ho�r'yIhMDs�L������4�~�AI��ʠX쳞 ���0��H�Ht��5gil����R_]W���,�WQ�Ɂ��#�&���c��X�@4ĕ]]�v0JѤ	[�=[�;�.�Är������(���0rD=�Q�r�6��W@���	�a�'q�y��A�����n�1��J�SA�I�%�	��黺q�s4����'|�A�1.u��j�eʖ�BdB}�r.���0��U���_�/�a����l�s��U�$k�6Ѯ�B>lo��K�UzB����+Ċ��HG�S*��-���2`�N%��R�l�Yib��tgż'�]U��07�!���K��?�,q־�/5�	<1��Lܩ7!܍ӬN#3_a�_�VJ&G�W�pm�A�v�;m"d�H����]糖�z��	KgC~����C~�V�'�]��W�z�@�of��E[����	��p/��Ik�;Fv�;������E��[��+���Gf�vS�������M��C1\�={�r��~D��O�5��l]���8<�������r{u��U��6�'G�?x(�b($g,��rUc;��]���~��6��e�9���U�hԈ)��	mPaT₩�-X�����S�'�I���Spv��8�_���C��}{���T��t�!����� ?�&4���5�>����\��-÷~�&������QK�Z�1i�˚��4���K]�D���A�D�|W�s��)����a�]Q��*&��ܿ*z�5	��U��@�'jM訪��r5i�$cm.w�m�X�P	�+k���R�j�Ѕ�o07 ��iH�4�����O��n�m�~�����g�I[���}�Q�}�N`�]2�!dch�ɺ&���Wy�WuP�+�ҷ��F�nRkIu�b�lߞE!�!��鶶�?�Qq�,�irS.�ܦZy�2F��~Tf���o�'���J�	�ś��l���uiP��FPJ�6O�QUf�/�G��s)�D/3�C��G�w;"=�e���kIx��l�	�%@�
���5Z���Em��&��4�l�:"(0_v}1���o��g�m�9c�(vH�y-I�p�F7��}Za�@AYOT?����ňxY=!�v&Z��}�e�������I�$��j��|p�j�)/o�-����>n�t�6~㾕�ً���`a	��n��߾?����^�Xč�\rVc0���L�W��4�h!���/���<nW�)�����x4ΥR��қ�ZQ�+�x���p����X��x!�lUˡ=^3���+
(�B!5s�B�!�����}�|�:�ƕD���������H����M�a�5���H�
p�L��4���=W˷��P��5Zb��*Ib���x�����m��JQ����EB�D-wK��@���՛��ТgC�yhN�p���"�Ik#<��y:	k1��]��V^8�m�=n��~���)!�b1�*!t� )|"+[4�VȀ�0(��k�Gť4\<�B]O%oN�b皥�H߈�5a�՞�O���w����a^�sAH�=���y ��F����!-(�n%Rn�q��FP	4\����հ�r���Y��`p���v{,���/���%2R&9|"O'u�y(�P̀��Z0{<頯��|�������Rd��P�݆�c��ո��W�u��*,�zFT6z���=8��Z����A?�����f6��1��Y����Q`��aD�Y$��*9��s�E%|���8}��zɒ�.F��ܳ.H���";i5��w����:y�0��������+��9s;YZ)���(�;�5�]z�JU���b�B3)���u�d;��҉�G�|������@� ��k'�Vp�&5���:����ä_v 2����ӗՄum]�v�x����W����*7e�ETr�7}F�*#m��N�r�zj8��n ���b�Y�OD4�����]c��ҏ�(����<j�ﴝ_4�螢���*��Oo�v�ka��%�p��� ���C3D�Ԫ��h�p����5]I1C�E�p�$�26~�GT&YR}���+J��X����������mk��HR�Oy��3[AP�	�1�\Usk�_[*��a" ž���由��oY�V�`h��6�Td	�ͯ�;���D���)��ߎ@������ct��.='��/�Ρ��/��!m�m�����k(��§��L��|�!�W�C	�";��_I�/�Ͼg��bȈu�����q'�v��uRa�+�h$Z�ԧ<�;!V��]ۼfE��e�jeE�qD󆃔Cr�Z���ĩX������Ee�h���ä�QY|ن^�P�e���Aೠ�-7P�,qf�¥�`�fӂWX�����&S�^/R�uJ�	��_WZ���-�zd�]k�DH�Ѷ.��W_wL�`��A~Z*�8ݧ��L��:��qT�|n�5\�޽�T�1�/�X����8�E|�5f1�n�kd�!ͨ�j*��{*D�Ki���eu�7�{�mzb/Gg���	��CQ-2�y�]�������>-7�U�78_ȗ��>Gb� =|��=]�CG��W�q�s��\߮�����2J�5�V�$v�(�1��T����ϖH�?���3,��-b��Ux)�L�SK�[j6[��<=��L���\R�z������"z�1��a��.��q-����� ������V�'⣝�mz�=�H����;�ߗ�D��=N��1����$�Iu�b
�s:盞��բ�D+��0E���m]��^<2�*��EL�oy�h�ұ��?� �����V���i%	9că��G	�Ѩw�q��u�"���a'X�X�6/j��.��n.��}�Rd0�+e[����̖d���X@uq���5M"gR���(���l"/ׅ�՚h���;\�0���A�uM�S�u�
n-K�7�ii��S��U��wѷv���r<buJx�wE����Ι����w�6X�8���zq{]��7w���R��1���̠[�|tU7\a�(��%���YKLT�XN�F�뻫��s�P���΍^�j�U$�x���V��l�q����`�e�_q�}^��|,�_���#��3�"���%}���6A�Ͱ��ƍ�^\�.	�H悰t���K��l�;"c��Z;�����\��r��Q�[6�w��-��D�杠��'��a�K_����%��u��VI��+��h���sN�~� ���s�'=��zH��Q�14��Yƾ��	�{ͣ��G`V�����x}0�	��&�R�~�;6l��U�hG��2L�[��[@sF\�ş�҅�����{~iϴg����(��y*���� ��d0�(��X\иݭ�qu��F|����\8�)����0��f�Ƒέ�?���$w��;��q�����šA��C�+������6H��_$w����<:�L46v�X�W����?I�{���t�q��.Y����)CMeJ�(�#f�5�a�+���B^*(!u������ؓ���-��St�� (�s��� (X��#��AyѾ���ږ�ˣ����p 'Hu��)Èdr6�7�V7�6*z����B����j+و�hmP@=�d��4�Y21+i���-���ULe�\<+\H:��}!pXΨ=������j�`��;>hn:?%�
8h�����h6�SM{�U}<�mzGʹ` g@T�ۯ�BV�d��qjj��۫&:�1��t��ôLv��?������:��NLU��ix�Z,늡+��t��J�Ϳj����j(*���A�	�L�X��%*,.�	WKϯ��X����MoM�;��������AD}j���ف��_���=)��>�TGg\.���A>�?��/��`�	o����~�e�͆=j�*.Ծ}u#�R��y��[H}��n�L^U�c.�j�䖭�?��$m(wq�*�;�z���&z|�i�j5F�a������|y��݉�X�XߧK<��c�6]4f
{���p��4�9|f�?:���&�$|�;��1�q$��e���c
�5�#��h�Q�)(�8#���^�[�M�e�'��acFD��N&�S��@���fC�'���U���ݪ���{}�)OYgP:X�˖Ft�%��ύ5[рf+�x(�"�ވA�q}jQtZ�:З�D���w�(�(z>���杏[��`�{�_�k���H̐�������qr���O���{=�
ˁ��"L�����]Gk�i �?1C��Lد�NԿQr�G����[hI�1K��&�%�;��9n�n�̓(޽��}�ڼ�B����a[���?�N^0��E�JK_]r]�4?%ܜȗ2��Ll����DN2)���&���V���d���,�\��f��
J��I��t���dE����U�q!OF�ӛ<y-P���:TK���o�U��qݡ}Z��~Y�)=�N��+��ɡ7Kñ���J�"��z�"��v{4q���]�Dz�<�n���yA��w��z���Ҡ=�[��U�<��%�e�N<�����l-�**t��1aL�Tzs�,ӽ�Ҳ� ��+����K�],��+� 6�I/��8��"Th{�h��JY���eSK	���b��@;�pW@!�P�Ǿ�J�i���|�Pѝ��~'��ϻ��z#M�*���A�~�BX�y�p"�kɪ�������L���Y}G#Pԝ;�i� �^{�D��s0-�ϊ��[��Ek�n�&h����}��-S���R�q#K�!��v@#*hϙ�R�8�����Ʉ�^YuNf��h"����}�m̿nhM/ A��e��e37���� �����y��}�6���5" F&��v�מ�v#���;S��XlxV16EB    fa00    1480��՜�A�IW��w�T�k9hEXd=��=Ŧ�2���XC�(z*�]���d����Z֙T�7Ɠ���[���*�d�RS��S�~��3?�sY�Ț2	1�xy�=�������ЂCPO���4L��<zI���ZvȄdο���ևt�E�Vuk}$x����Ȑ�*:��M�9��`������Z�b�p)7���\E�aC��}�M:���cq�3}<������L����[!6��
�]D����3s��q�)L�k��}q�
N҇���Zh���M���ѩ�;�W��qyFZU�1��������gB��������fM<��.�x�z��t�Z5Y�\��c�z]9���+75>сߥ3��&��G�iKh"�>�oq���|Yk>̏)�Ϭїhr�|"!6pn��/;
�}������!"��'��~H�ۦ�$~n�6X�C��6��zR���OR9�c�ݗx,�`�N�!�%�PբlOkY��%�����������ό$���8d��L�
 �(D��_Ĥ0{ס�;k9�8�O�.4s��FldUK��'��q�f�zj�0��m�\w'�c��]հ�Ⱦb�z��M�<��9�s����m�@��L� ښ��_��ݹ?�
����x7�O��|k��`���!��W�:P8���o��*�A˞���|��=+��f���j�Lٓ��{gY{�C�^� !���{h��Q����� 1���@,YL�Zo,:����/��	XP9pZ��9�
)j��Hu���!�'���q�@+�rm]�1nk��8�x�Mp��.-E2��w���?@��VZ ���P���+W���;m#�O���3�3Cd���R.[�J0���q�=����4e��ٜ��ca���D�$S��y��ŅYDn��-�4U�ڱd� "�����7���rR+�ѫ��s� �|����E^�Z���Rx��e������eX�FG5�>Qj�{�?�I5�c6�T���*	"ۈ�@�XN�� ��J���'�q���\�9"ä�͘&@��7��:e� 0��F�R��^�APAm�TB��F�K6�¤Ef.ⶖ~�_
����B��;Qf���D��ʜ�,�N�ȉ��e�(�Tl��(�L������?9�Ct�:T}���ę���5�T�*��N���$�<�7Z������1��D�CC^��n�pǃw�(=�6%��Y�ů,��=Q�W;� ��,�3#�$�՝bQZE�j��ﾧ?JC��C�º%E�H��{K�8$��o�ۆ��h�3F�A�2���l��`���o�G�t�k8����f���ϓW9%W���5-2��/Ѓ�֮8K�����L�6�`���څݾ��&��A� R�Ԓ�i�Dx������.4 ��`�y������"m���y�.q�a*}���5q��/��נ�wx�M��WII�W!�Mb&�tT��=U	4y?��c�0�b��b�$�T�{��C�+��*�������d���ɳ�g�F� ���p	u�����_q"����V�2����;j ��k��]���w�v.e��%J�|;8�	$� ���=*w1�YS�B�_�4V�����*d�hh�U��c�u�~̭���v�+K8����	π� L�G[��ܸ#_������;���� �M������<�λ0��%���_~�	������v an��#Y��쐑��g+�.1��rX�A�vg<����=��>�7�z2��B���yC+d��5<� �3�tC�?�C��H�P����x'ރ��mg\�H��uu��]�ߴ?�!0~�t[��AE�QW�8�l�4{��G��3?�ܵH0���~q�Y�%#K�:ػ�������l�_ɂ���vI�J�)5T']W�@8�B�b��<A )q���a9��D��'��z���P$���e7�ѻ���
�1^����Rhj��ٗBb�	IE�Y��2Hҽ�� >��q9��kTc�C����2D���r^���{?g�|u�9c��ZE�(�Z)2��u���2�F�~�r|UTq�A� �`�ؓ�y��j��1��\�z]}�*"ܙ l�cG�%����r|<^hO>:�D�"N�����FYe8���H��R��h�7@����X��f�o����?<LFO�W!�2V�T��T��J ��ZE����d��B%���f��Y��C�v�dʗ�:D ��(2?�|����j��om��p��,'H�9gP��	�w@��h3͹:��X�C���W��|�r嚂o� Ղ /J�{���ů��3'k�V���'*��i�O���V5�h�4�W2��Y�4��U���(c�m�>�-^O�y�4Zv�b�K�� ��4	ClO�XX��8�F7!w}$^�T�E�@@\�a�P0�a�W����"�`�X~��f��
h����ܩ"^��i,��B�3��,�9��mqy�3��dz;�mũ���W�k��;��N��k��@WvHq��-����|�Bէ3�{&��Pm��RF�&���#���,�*K����RfJC^a32��HIW��3�^��:�����)ҿmo\!�����8ΐxF��O�'gyB-�ͩ�d�t�]����g�j�c�&Ow�`���}��&�}J�>�D϶Wp|�a�퇖۞��iJ�#ĉ\����6�H�#����d��3K�%R�����'��^�*��az����7���W7�2��V��qfc�8�Eʴ���eK��Y�
H\�w��Q`�uf��J^r99��Jʊ�"s�j2-���0l���!B�A;���� oi@S_l�h���c�k�IŁ�A��5#�PB��Ĳ����#����\���!Ô�c����=}����4�~1K��~pi��$
����� ��O�vi�=\?�։|���31��e�������s�j7���u�
. w�8��%���y	���<���ɏ�ذi�-��C# �L��nF�v�k픖������ޠJt��~��,"�U�V��^���Q}x�(uw�(����X�PZ�ID&<Є��&C�q���2��]���u�A�AQv��BAX
������KM&C�=x�I�O�O)���\��_9�}g\�WV>��./C���,]�"'��B��H�sD��9ӵ����רAa��X؜r�^z�_4'����G���F�;G���W�\�)��Mޜ��Y�5}�.�iH�D�c=5���Q�"1�?���Ν�XK���K!�VWe�[L��W��3��i�xH4ב���hI����q6�>1�w�N?q1g;,TxzP�p1W:歄�g�U������)�+ܷw9�Bّ��!fc�"ݲ}��Y�`6��wSv�C��r.̘������^Ҋ�~c\���ej�p W�Y��n�L���5���w xR������CHq�G��WJăŢCO~X ��V�K���s��Ѷ�Ls��M;�g�,��Q��h(u։ 8���vn]�� ���9fp�� �@r�~��D����r���q��$��r�F	�Ոܼ�*�N�i⣿�,Q�D!3..����䜿��*�.�F��JrO��9�uy�QC�%�n�d��*/���1�6���Vwތ�1���=���芃}�ayv-:@
���ET2�i�᣹���;��~�sv�զ¨���R|$�ϙ��Ƌ~�N�b��:I��s�u�+�����]4����@���W��?����L4Uɐ����^H>Eg�Q�-�)g�1nl�`ƹ7a��=7�~��O�����w�5�0?OV$`K�Z�x}>��������]��(�1]Ӳ܏&iNܸڸXTX��4����=Ρ��S#��"&nC}9@L�o!�)@��f�������B�ƾi��b�,�?z]�o8V�X�!�نU |����t�W޶H'С�J�Y2H`(Y�Ó��@fd5 q�\�H���W�Bl��^�2Et�01�?�i��y՝���2��wk�=�n�u�y!Gz��ע�gѰ&;2#�+M1�næž�$,I�E�t����6Ć:gAG<{;�_'6��;Ș�G@�'�	��\\�(��=���n�*%K�A'@��ox�<ԣf�0#[��~��xԑ�0ج._֬/����� ^u;�XM�A>����U�J�O.JӞ�ꢪ�k2�㰢(�j0t9<����>�,�R�Z���T��^6�>�h]\��zh	˙e!��o��$
)ѼE����A��"S�Ƒ$��9����cS��x8Ml�7:Q�e�ZW z���܁�UZ�?�WX�Բ�L�wyrr6�+�\[`|h=/�[���nj
i��|p��LT���������Җ���%0�g�G��J\�'�}Y�~t���$2D1��d�
K�Ǘ�Z>�i��kU7?�_(p+Ee�O���Jt���(���>����TY)���j�&�J�*(���@D�_rS4�Q����w�*�5Xmd:�	(:�D�S�ADyYd|<	�Z�b�M�Z_`���Q����֭�YVUq>Hd{�O]btxjױ_;0j��![��L��B!�����.i����i��?�Șw��[���G>��}��A��gV�k��A|4���=K8�����!m"\�C�ZQ�J�y���l�l �"6!-���\�]Y@�s���x�t1ӱ�g����FCv���b|w<oL���(���Ö��t�r"��%Nb���1�8-����x�}�9�x\���P�vu>_����4�֪֛\F.mI^e�&X��gH@��S�~Zͨ����6��E-"�hT�jvQ�a���v�E@R��(plˌk�3�of��;L�b[w,г/T?lq�}���P ��:��=���Ễ�Rh��� iW�$�y�ׇF9D�?q�$"0�E�	yDs�j��`ʓ�跶�S�Y��f&챸�A��	72�nx#K��m���+~��r��Hl^g-Ђ;�)��n�Bb�cl���	�T3O�Q
<\�b��A���fAblY�`ʢx���΋��0F�Q�*�Zq˹���聥`6Jz�MJ鿈n|��_��ծ������P����+ �)p��V� �!�<��U�x�\T��}��;ǐ�9�ٰ��R��^:o�2���i�ψ���[/ڧ$��mիJ+��jXlxV16EB    fa00     d50ȋ�`��a�AkG2C�&j�
M�����d1���c�^�Ǯ Xh����L/��E �'�_G�L%7��Yt�:g�\h��8H�ֵ�N���7�^%=������o"vSZ^�);Ѳp8�Ԕcڗ�?�[lII�/�f9���c��ԛ�/�
�ʍđ	ϖ�JW)�ǉm���=0a����WP56��2�Q��I<z?\!��=:��;v��qIq�h�|9qeC,��9�z觠�'��]d��Kc2�y�)܎Q�/PJ�D>yKC)Z���=<�Id�ci�̜��U�5/�>.��8<4��Ą�-X�=$F��E@��o-�l�V���V�/�|�8�/������6Sf�����H�0�"Te^O�J�}�>7$U��_�0��▝��yk&�6^�`D�x�Ċ�K�r`�D_���FQ:Rd}kH���	8��).��U<�fq�as�)R�#M|�;��K��l4���攒��K�B3�,ѥ������c�@i��3�|Q�s��U����b�p�o�_� ��zCM|S'��)ER�ʓ8u��H�O<KNΕ���]�Ċ�L�B�2���e�v=2�%O����ܠ"޸H��q��ҥ,����eS�d;{�ze?C	@ؓ����$R6���&���r�W�*�Eg��r
���(�3*8�t(�V���� @t�w��'o-�d�Bj�"�g}�(Y�v���W�X�{���{G�,��{(���r�ހ2a���k��L�\�k5����N1s�a�6H��-�Uf'��n޲�^��.�*&깑m>E���4��\4��ݬq�X�����*n#N�۝8�^��3�,���	#˧���,�&T�W��HX�Z��5p9�ܔwp��&�Jb3#�1���W'�NkZ��f��D�W�֜{�W����/:��y���N��w�׋Kw�6ח�{�檎5�\f3#\a�d�2���;���bV>+��Z�=��P8��>�Z��N��Z7���n?�Xq�� h�Q������E5	R�4|n D�>�&=qz
Q¤^fx��C�Z��}�U�EJq���p\�� �¥t��k�������T	�)�	.BW�b|��BOP^��U����OÞ����;Ǣ"�J���b���6�I��:��[]�/<�
D�9�B��� 6��:���؂i�*,��9�m�Z�0 6����)}�5��;,o^���'�E>R���8\%�dDX�%��T�_�!�8܄S4b#1�+�] �[��t��޳Ɩqxu�{�m�fɧ;B�};�����_��.�w�
#ƨhuK���N2dḧ؍�<	t�$@�S��B��a|ˀ���Ѵ�dJ6g��� .mI=��l�o����e���-q��*�\�	������$Yٓ�X�*���W��7��&���tۙ��qLf�J�˛��Lf;�|� ;Q��I�-aj*��t�	zr~�:�6i�!� H��Lg�!���ՋÓw�����}%�d��n��5~M�'�p�����a�J_�#��
o�B6LE��_��x(��WT+~�l-�6� �mH>�/}*��Qʿ88[~�w�2 �[�TlbUt<�e,s>:?�[��f����o
��H�z>A��NgI���hW�P���@���������GܳL^��uL|�"d�Z;�լ�N�s$N�)�(��$Ͻ��2&qvC/a��ي�h��E#*�L�I�3�ߴZ��[P#Ph-�^qa:'���^2��1��I�aU��BG�{��,�>[�rgs�w�U����F��.z����N��8�S^�;m�#����V�A���e��Kv�.b#��
�v��:~ӛx��P|P��.{4ĩ��_B-Q'�;���\��-�eZ���\�Nv�|9�)��c?[���󦎩���MG%��
���E-T�q.���]/�ڏ�X%��g���#bB��>�G�v� ����h��5O��j�6�P��1r��F�H��%z�N|����3/g�+���r���w�����
��9t�4���$�����GX$~&���e���/Z�w�.hv��l�%2]��B1�,���U��0�x��ٸ&U)��8�C!�2��Nے'-'����Q��=|��A\.�F�G�k>��s�m����j;k�{�;�	h�Ɵ�A���q��U��-uI[���]�R=�W���;�KX�S�=�*bl�L�LaD	�J��16�� �_O�������J�#\�63؃oԊeｶ` ��������RSW�τc�)�
�RI���;�����f�|��U�X�����v�J��G^p�R\��'׹��W�@0��pZj�5<N*�gaLot��:��n��=��X:�B��I�xq��_��_�;�BH�x�/�9�����(� ����7��Y�i��)E>��e����c�� _����[��w$�KP�bMhny���ិ=�c����S�QEQ�ߊH\�<���@a5��EJ1�
�0gؿM����Z���IL�-�p24�J�~7f��J�❹Hi|���_�2��-�t��oñ����2{���S=���
BO�>��!�&�c.��Lϒ���J���|�o\0����޳xQl^�0`>i9'X�l���FO�B
�ܔ� ���
s`kr�X��i���)��OV�iSDz�CU��(<5�-�Pcߠ}D����D<N���?^�1��wڙ�t?M@K�~4Y��F�*EU$*]��<Sn$�l����D��\��3l��m�MXkH D�|��"J>0D�7WN����[�P������Z��uBޤ=��S�-����)�.a�K�v��$��Ar0,IdKy3Ɗ�V'����+�6�*�H���'����?��&1��o��/�>��ߢ%�6�r�X��^0�N����Ī�foƘ���¾�/��)�� �N}�7��f�w][JY�$���޴��O��V����a�8�x���!��BU�Qo;ӷ*ލ�3�D�����������i�4�~�*�S�i|��@�E�5��Жs�Ğ�IԷV��ŔDC�+b{�H�u���PuC'l���i>�R�]��X�aVM��~�h��Jj�����EgF��זO��@?���� �x!K�2�e�F0�ѵ�25ꝫk���7�*�O�fKz��k�A}��r'-�Iჴ�=�/�s�v5\
=��/��{-L~Lu�f��Jj���Q�|�u� =ݩB�_�r9�#_�tC��vRȉ͖.L�)xw�����7��ҵ[)5kB$�z���%wV��K���(�n�w����$ń�F��/Ŷۈ[�k����j���^L�fb�&�z�u��XlxV16EB    9230     c80a@]��|������a{l6�R�O��v0a��#���|D��+�K/o���\�|��]�i�h�*	J��X����h&�:S[?#_���%i��^��[����������\�=蔒�
��ӥ\%ʯ���bv+�q�R��/aM���Y��6*�(g�Mv���*p%��a	fC�p��7q�O�^r��N�"�^��V�O�4��rTB�Eل!���;�s��*,�'8r�-;_`Ò0K����� ���JC�I��P���s��Ĺ�/x�\��O�>��"M%l3���Q6��i�*�U��4ÑD��@p����)��7��O����i�E����ş�G��*�����N�A�7ن��v���@����i#����!S�>Ȥ��=GZՒi�:��#��+AQu�|ݕ���n5���I���J��Ot1ᷣFk�����Ã�͂dk�%�|��G�>�&j�2X��}1��=���|��ҹj(r�i�q�	,R�y�:H'��2��غ� 0�XZm�>��.�SW@߈��H��XE�Φr�F��يⶍ�������U��� j��a_�k�̍�5��`[��3��!�Sx�����]n���p�.���'�;G�A��R ��[H�j�Q�6���*k�Xr�v��Gú;�"���\Y�>��҆�:b�K�@i?t� <O��#��W�^���7b����}����dn<�jB�y��H���c�ܶkĿ]!(~=����(;	����U���\�"����p鑿M.k{�JR�A-�\~�Dc�)i�N�Kq8=�I�*Niz�u���쿢
��%	N��%�8��`W��
�����bI�3��� B�^��_B��P������Μ��{z�.�tQbo��q@���Ŗu�h������w�* :�]��y�G�$6�5[�X��ת84~�o��>�;iG��E�=`�����tj�C,r1p�U+�����I��w?�\0�>"遽=�]�+�`��.=��d��b�(�z�o�X	��T��?|[�p�Ǘy�$R$�}�]F�#���n
x�1�=.o;�in7�18�;[UEsNJ�v�:�GG�ֱh[�����ך2I���,&�y➝l=�и�G@�� }_=�}�q�Cjw:�.|T*�`��N��) Gal�ff9��a=���:��c�'�͍��s�0\v��$�� �5����1 ����,�q^z���!f4&{S����!��
2������G�ܻ#�%����&8� �kT8�|�qI-��\��m�� ��	���ŵ���B�&L���f���◘��t�n㥺�<����{BYz��R��4B��G�|�����d�����1����[;�(K*{/�{�MO���B,����1��V~�c��U�dV�'��Ɣ3*̔�N�Ȁ4El�K�lpP39�AR$l3r����&t���<,B.�H@M��M(�/���)�va���pȝ��8ց� O'������_$�x�8��-��7L�3��gxo���J�����	6�?/̩%ϣ�n���<|8G2=�g�^{�f�)`,~c�->�0���U��K)��~�%�W[���1�I���o�^����V�j4�3��~A�G��p;����MR2��]����Fݟ�aj���D��z[��4�$�a�.[���a�&�o?�d���)�K�G���V�J@��/6O��g�Kʛ!0��@\D(0Td�I.��&��sp6Gˏ�E������8ՠ*pfc�2<��[�4�R����L��9$w~ֱ%��*�JP�unx�?'?�)��^�n\� =�Ưn M h֛�|�j��C �d��+��o�Qm��?��*F_U<��d��m� �Tѻ�q�kU��
`�������i,V��Ti�_�����f#�l�%��nW��I��	(�i��A� wJ�5�[��m��)�ޑf-j< ")��ǉ�p���,ƛe�b��M��L֙	 "�r@�j���ܧ��3�2⋊	. :=�Y;>R�3��[�7t�^���'��O�8�g��
%Xx��sb�Ղ��]��˭d�Bd�������א��*��Ջ��BBrt<?�g(��\msaJ��3b�|� �9�s4������,�Z��^����Z�)��� N����$��cJ^��ؑ�U~�2�DD����tYÈ/<��O�'�Z�oyny���'qKϿX�$�p٫`�f��m��Ԥ���[�j6������&}�+��{��.�tG�i��9];ݾ���F&�~�d�D9�b�f�}x�Xg6[n�G�1�1�'��@�����À*3��c[Kv&R����$�|�S��l}��녚�@1�(�5j�=W��T��Dp@�񁑐��#A��4F��S�M!/�7��m�/{�f
p���E�?mT)��G�6��q��<'I�I�{�g������:
F��Q�!�ñ��T�R��~/e.ށ�(�?��{���~ȞnU�&�M�$�-O�2������ά�ӃU��<7�Z2��h[?$=�b�}�c�U�������2�@�Y�>J(�^�Jj�;���Ch���9+�&�< �*�'��S���P2�`N�T���i��)T�d�1������	�S7j�������L�Th�<�O׷�]@�=| ��tB�;mV��X�� ԤYV��\���BX���f��@�ӳ+2���֫Y-���W~/��
��Y�_���4�ql���V�/���N�J�X[�0�׻�(�� ��^��x����P��]h<�aI3Im����9���a�Td�P�K�͂s�IL ��u��^rYE{���&��i:ZKEs��ykZ�PV"N�t�����O!0p�_:j f�Z�2�Q8��9���2����6Ur���i�$O��2>�ilD�^�����2%��I ę|%�C�"F<��1��-��R�y�-�g�C?nr09s�X�t�Y!��cuR�kI���lm¡�Z�In��\;�E�ě�{�-���U�:Iб%��>N��<,�6r��T�\/τal~5�R>���Q���5N5���N�}��+�[��&{���Ȋ��11π�Ax[$������	�{0���[�C�=x�+5��>���ʒ9��
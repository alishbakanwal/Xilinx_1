<<<<<<< HEAD
version https://git-lfs.github.com/spec/v1
oid sha256:47490f68635ee86f6f2cc94846f2153b829d49e8db82c5bfe344f2362031c842
size 92662
=======
------------------------------------------------------------------------
--
-- Copyright 1996 by IEEE. All rights reserved.
--
-- This source file is an essential part of IEEE Std 1076.2-1996, IEEE Standard 
-- VHDL Mathematical Packages. This source file may not be copied, sold, or 
-- included with software that is sold without written permission from the IEEE
-- Standards Department. This source file may be used to implement this standard 
-- and may be distributed in compiled form in any manner so long as the 
-- compiled form does not allow direct decompilation of the original source file.
-- This source file may be copied for individual use between licensed users. 
-- This source file is provided on an AS IS basis. The IEEE disclaims ANY 
-- WARRANTY EXPRESS OR IMPLIED INCLUDING ANY WARRANTY OF MERCHANTABILITY 
-- AND FITNESS FOR USE FOR A PARTICULAR PURPOSE. The user of the source 
-- file shall indemnify and hold IEEE harmless from any damages or liability 
-- arising out of the use thereof.
--
-- Title:       Standard VHDL Mathematical Packages (IEEE Std 1076.2-1996,
--              MATH_COMPLEX)
--
-- Library:     This package shall be compiled into a library
--              symbolically named IEEE.
--
-- Developers:  IEEE DASC VHDL Mathematical Packages Working Group
--
-- Purpose:     This package defines a standard for designers to use in
--              describing VHDL models that make use of common COMPLEX
--              constants and common COMPLEX mathematical functions and
--              operators.
--
-- Limitation:  The values generated by the functions in this package may
--              vary from platform to platform, and the precision of results
--              is only guaranteed to be the minimum required by IEEE Std 1076-
--              1993.
--
-- Notes:
--              No declarations or definitions shall be included in, or
--              excluded from, this package.
--              The "package declaration" defines the types, subtypes, and
--              declarations of MATH_COMPLEX.
--              The standard mathematical definition and conventional meaning
--              of the mathematical functions that are part of this standard
--              represent the formal semantics of the implementation of the
--              MATH_COMPLEX package declaration.  The purpose of the
--              MATH_COMPLEX package body is to provide a guideline for
--              implementations to verify their implementation of MATH_COMPLEX.
--              Tool developers may choose to implement the package body in
--              the most efficient manner available to them.
--
-- -----------------------------------------------------------------------------
-- Version    : 1.5
-- Date       : 24 July 1996
-- -----------------------------------------------------------------------------
library IEEE;
use IEEE.MATH_REAL.all;
package MATH_COMPLEX is
    constant CopyRightNotice: STRING
      := "Copyright 1996 IEEE. All rights reserved.";

    --
    -- Type Definitions
    --
    type COMPLEX is
        record
                RE: REAL;        -- Real part
                IM: REAL;        -- Imaginary part
        end record;

    subtype POSITIVE_REAL is REAL range 0.0 to REAL'HIGH;

    subtype PRINCIPAL_VALUE is REAL range -MATH_PI to MATH_PI;

    type COMPLEX_POLAR is
        record
                MAG: POSITIVE_REAL;    -- Magnitude
                ARG: PRINCIPAL_VALUE;  -- Angle in radians; -MATH_PI is illegal
        end record;

    --
    -- Constant Definitions
    --
    constant  MATH_CBASE_1: COMPLEX := COMPLEX'(1.0, 0.0);
    constant  MATH_CBASE_J: COMPLEX := COMPLEX'(0.0, 1.0);
    constant  MATH_CZERO: COMPLEX := COMPLEX'(0.0, 0.0);


    --
    -- Overloaded equality and inequality operators for COMPLEX_POLAR
    -- (equality and inequality operators for COMPLEX are predefined)
    --

    function "=" ( L: in COMPLEX_POLAR;  R: in COMPLEX_POLAR ) return BOOLEAN;
        -- Purpose:
        --         Returns TRUE if L is equal to R and returns FALSE otherwise
        -- Special values:
        --         COMPLEX_POLAR'(0.0, X) = COMPLEX_POLAR'(0.0, Y) returns TRUE
        --         regardless of the value of X and Y.
        -- Domain:
        --         L in COMPLEX_POLAR and L.ARG /= -MATH_PI
        --         R in COMPLEX_POLAR and R.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if L.ARG = -MATH_PI
        --         Error if R.ARG = -MATH_PI
        -- Range:
        --         "="(L,R) is either TRUE or FALSE
        -- Notes:
        --         None

    function "/=" ( L: in COMPLEX_POLAR;  R: in COMPLEX_POLAR ) return BOOLEAN;
        -- Purpose:
        --         Returns TRUE if L is not equal to R and returns FALSE
        --         otherwise
        -- Special values:
        --         COMPLEX_POLAR'(0.0, X) /= COMPLEX_POLAR'(0.0, Y) returns
        --         FALSE regardless of the value of X and Y.
        -- Domain:
        --         L in COMPLEX_POLAR and L.ARG /= -MATH_PI
        --         R in COMPLEX_POLAR and R.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if L.ARG = -MATH_PI
        --         Error if R.ARG = -MATH_PI
        -- Range:
        --         "/="(L,R) is either TRUE or FALSE
        -- Notes:
        --         None

    --
    -- Function Declarations
    --
    function CMPLX(X: in REAL;  Y: in REAL:= 0.0 ) return COMPLEX;
        -- Purpose:
        --         Returns COMPLEX number X + iY
        -- Special values:
        --         None
        -- Domain:
        --         X in REAL
        --         Y in REAL
        -- Error conditions:
        --         None
        -- Range:
        --         CMPLX(X,Y) is mathematically unbounded
        -- Notes:
        --         None

    function GET_PRINCIPAL_VALUE(X: in REAL ) return PRINCIPAL_VALUE;
        -- Purpose:
        --         Returns principal value of angle X; X in radians
        -- Special values:
        --         None
        -- Domain:
        --         X in REAL
        -- Error conditions:
        --         None
        -- Range:
        --         -MATH_PI < GET_PRINCIPAL_VALUE(X) <= MATH_PI
        -- Notes:
        --         None

    function COMPLEX_TO_POLAR(Z: in COMPLEX ) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns principal value COMPLEX_POLAR of Z
        -- Special values:
        --         COMPLEX_TO_POLAR(MATH_CZERO) = COMPLEX_POLAR'(0.0, 0.0)
        --         COMPLEX_TO_POLAR(Z) = COMPLEX_POLAR'(ABS(Z.IM),
        --                              SIGN(Z.IM)*MATH_PI_OVER_2) if Z.RE = 0.0
        -- Domain:
        --         Z in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function POLAR_TO_COMPLEX(Z: in COMPLEX_POLAR ) return COMPLEX;
        -- Purpose:
        --         Returns COMPLEX value of Z
        -- Special values:
        --         None
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        -- Range:
        --         POLAR_TO_COMPLEX(Z) is mathematically unbounded
        -- Notes:
        --         None

    function "ABS"(Z: in COMPLEX ) return POSITIVE_REAL;
        -- Purpose:
        --         Returns absolute value (magnitude) of Z
        -- Special values:
        --         None
        -- Domain:
        --         Z in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         ABS(Z) is mathematically unbounded
        -- Notes:
        --         ABS(Z) = SQRT(Z.RE*Z.RE + Z.IM*Z.IM)

    function "ABS"(Z: in COMPLEX_POLAR ) return POSITIVE_REAL;
        -- Purpose:
        --         Returns absolute value (magnitude) of Z
        -- Special values:
        --         None
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        -- Range:
        --         ABS(Z) >= 0.0
        -- Notes:
        --         ABS(Z) = Z.MAG

    function ARG(Z: in COMPLEX ) return PRINCIPAL_VALUE;
        -- Purpose:
        --         Returns argument (angle) in radians of the principal
        --         value of Z
        -- Special values:
        --         ARG(Z) = 0.0 if Z.RE >= 0.0 and Z.IM = 0.0
        --         ARG(Z) = SIGN(Z.IM)*MATH_PI_OVER_2 if Z.RE = 0.0
        --         ARG(Z) = MATH_PI if Z.RE < 0.0        and Z.IM = 0.0
        -- Domain:
        --         Z in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         -MATH_PI < ARG(Z) <= MATH_PI
        -- Notes:
        --         ARG(Z) = ARCTAN(Z.IM, Z.RE)

    function ARG(Z: in COMPLEX_POLAR ) return PRINCIPAL_VALUE;
        -- Purpose:
        --         Returns argument (angle) in radians of the principal
        --         value of Z
        -- Special values:
        --         None
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        -- Range:
        --         -MATH_PI < ARG(Z) <= MATH_PI
        -- Notes:
        --         ARG(Z) = Z.ARG


    function "-" (Z: in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns unary minus of Z
        -- Special values:
        --         None
        -- Domain:
        --         Z in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         "-"(Z) is mathematically unbounded
        -- Notes:
        --         Returns -x -jy for Z= x + jy

    function "-" (Z: in COMPLEX_POLAR ) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns principal value of unary minus of Z
        -- Special values:
        --         "-"(Z) = COMPLEX_POLAR'(Z.MAG, MATH_PI) if Z.ARG = 0.0
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         Returns COMPLEX_POLAR'(Z.MAG, Z.ARG - SIGN(Z.ARG)*MATH_PI) if
        --                Z.ARG /= 0.0

    function CONJ (Z: in COMPLEX) return COMPLEX;
        -- Purpose:
        --         Returns complex conjugate of Z
        -- Special values:
        --         None
        -- Domain:
        --         Z in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         CONJ(Z) is mathematically unbounded
        -- Notes:
        --         Returns x -jy for Z= x + jy

    function CONJ (Z: in COMPLEX_POLAR) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns principal value of complex conjugate of Z
        -- Special values:
        --         CONJ(Z) = COMPLEX_POLAR'(Z.MAG, MATH_PI) if Z.ARG = MATH_PI
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         Returns COMPLEX_POLAR'(Z.MAG, -Z.ARG) if Z.ARG /= MATH_PI

    function SQRT(Z: in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns square root of Z with positive real part
        --         or, if the real part is zero, the one with nonnegative
        --         imaginary part
        -- Special values:
        --         SQRT(MATH_CZERO) = MATH_CZERO
        -- Domain:
        --         Z in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         SQRT(Z) is mathematically unbounded
        -- Notes:
        --         None

    function SQRT(Z: in COMPLEX_POLAR ) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns square root of Z with positive real part
        --         or, if the real part is zero, the one with nonnegative
        --         imaginary part
        -- Special values:
        --         SQRT(Z) = COMPLEX_POLAR'(0.0, 0.0) if Z.MAG = 0.0
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function EXP(Z: in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns exponential of Z
        -- Special values:
        --         EXP(MATH_CZERO) = MATH_CBASE_1
        --         EXP(Z) = -MATH_CBASE_1 if Z.RE = 0.0 and ABS(Z.IM) = MATH_PI
        --         EXP(Z) = SIGN(Z.IM)*MATH_CBASE_J if Z.RE = 0.0 and
        --                                          ABS(Z.IM) =  MATH_PI_OVER_2
        -- Domain:
        --         Z in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         EXP(Z) is mathematically unbounded
        -- Notes:
        --         None



    function EXP(Z: in COMPLEX_POLAR ) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns principal value of exponential of Z
        -- Special values:
        --         EXP(Z) = COMPLEX_POLAR'(1.0, 0.0) if Z.MAG =0.0 and
        --                                                        Z.ARG = 0.0
        --         EXP(Z) = COMPLEX_POLAR'(1.0, MATH_PI) if Z.MAG = MATH_PI and
        --                                        ABS(Z.ARG) = MATH_PI_OVER_2
        --         EXP(Z) = COMPLEX_POLAR'(1.0, MATH_PI_OVER_2) if
        --                                        Z.MAG = MATH_PI_OVER_2 and
        --                                        Z.ARG = MATH_PI_OVER_2
        --         EXP(Z) = COMPLEX_POLAR'(1.0, -MATH_PI_OVER_2) if
        --                                        Z.MAG = MATH_PI_OVER_2 and
        --                                        Z.ARG = -MATH_PI_OVER_2
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function LOG(Z: in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns natural logarithm of Z
        -- Special values:
        --         LOG(MATH_CBASE_1) = MATH_CZERO
        --         LOG(-MATH_CBASE_1) = COMPLEX'(0.0, MATH_PI)
        --         LOG(MATH_CBASE_J) = COMPLEX'(0.0, MATH_PI_OVER_2)
        --         LOG(-MATH_CBASE_J) = COMPLEX'(0.0, -MATH_PI_OVER_2)
        --         LOG(Z) = MATH_CBASE_1 if Z = COMPLEX'(MATH_E, 0.0)
        -- Domain:
        --         Z in COMPLEX and ABS(Z) /= 0.0
        -- Error conditions:
        --         Error if ABS(Z) = 0.0
        -- Range:
        --         LOG(Z) is mathematically unbounded
        -- Notes:
        --         None

    function LOG2(Z: in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns logarithm base 2 of Z
        -- Special values:
        --         LOG2(MATH_CBASE_1) = MATH_CZERO
        --         LOG2(Z) = MATH_CBASE_1 if Z = COMPLEX'(2.0, 0.0)
        -- Domain:
        --         Z in COMPLEX and ABS(Z) /= 0.0
        -- Error conditions:
        --         Error if ABS(Z) = 0.0
        -- Range:
        --         LOG2(Z) is mathematically unbounded
        -- Notes:
        --         None

    function LOG10(Z: in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns logarithm base 10 of Z
        -- Special values:
        --         LOG10(MATH_CBASE_1) = MATH_CZERO
        --         LOG10(Z) = MATH_CBASE_1 if Z = COMPLEX'(10.0, 0.0)
        -- Domain:
        --         Z in COMPLEX and ABS(Z) /= 0.0
        -- Error conditions:
        --         Error if ABS(Z) = 0.0
        -- Range:
        --         LOG10(Z) is mathematically unbounded
        -- Notes:
        --         None

    function LOG(Z: in COMPLEX_POLAR ) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns principal value of natural logarithm of Z
        -- Special values:
        --         LOG(Z) = COMPLEX_POLAR'(0.0, 0.0) if Z.MAG = 1.0 and
        --                                             Z.ARG = 0.0
        --         LOG(Z) = COMPLEX_POLAR'(MATH_PI, MATH_PI_OVER_2) if
        --                              Z.MAG = 1.0 and Z.ARG = MATH_PI
        --         LOG(Z) = COMPLEX_POLAR'(MATH_PI_OVER_2, MATH_PI_OVER_2) if
        --                              Z.MAG = 1.0 and  Z.ARG = MATH_PI_OVER_2
        --         LOG(Z) = COMPLEX_POLAR'(MATH_PI_OVER_2, -MATH_PI_OVER_2) if
        --                              Z.MAG = 1.0 and  Z.ARG = -MATH_PI_OVER_2
        --         LOG(Z) = COMPLEX_POLAR'(1.0, 0.0) if Z.MAG = MATH_E and
        --                                             Z.ARG = 0.0
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        --         Z.MAG /= 0.0
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        --         Error if Z.MAG = 0.0
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function LOG2(Z: in COMPLEX_POLAR ) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns principal value of logarithm base 2 of Z
        -- Special values:
        --         LOG2(Z) = COMPLEX_POLAR'(0.0, 0.0) if Z.MAG = 1.0 and
        --                                              Z.ARG = 0.0
        --         LOG2(Z) = COMPLEX_POLAR'(1.0, 0.0) if Z.MAG = 2.0 and
        --                                             Z.ARG = 0.0
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        --         Z.MAG /= 0.0
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        --         Error if Z.MAG = 0.0
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --        None

    function LOG10(Z: in COMPLEX_POLAR ) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns principal value of logarithm base 10 of Z
        -- Special values:
        --         LOG10(Z) = COMPLEX_POLAR'(0.0, 0.0) if Z.MAG = 1.0 and
        --                                               Z.ARG = 0.0
        --         LOG10(Z) = COMPLEX_POLAR'(1.0, 0.0) if Z.MAG = 10.0 and
        --                                               Z.ARG = 0.0
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        --         Z.MAG /= 0.0
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        --         Error if Z.MAG = 0.0
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function LOG(Z: in COMPLEX; BASE: in REAL) return COMPLEX;
        -- Purpose:
        --         Returns logarithm base BASE of Z
        -- Special values:
        --         LOG(MATH_CBASE_1, BASE) = MATH_CZERO
        --         LOG(Z,BASE) = MATH_CBASE_1 if Z = COMPLEX'(BASE, 0.0)
        -- Domain:
        --         Z in COMPLEX and ABS(Z) /= 0.0
        --         BASE > 0.0
        --         BASE /= 1.0
        -- Error conditions:
        --         Error if ABS(Z) = 0.0
        --         Error if BASE <= 0.0
        --         Error if BASE = 1.0
        -- Range:
        --         LOG(Z,BASE) is mathematically unbounded
        -- Notes:
        --         None

    function LOG(Z: in COMPLEX_POLAR; BASE: in REAL ) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns principal value of logarithm base BASE of Z
        -- Special values:
        --         LOG(Z, BASE) = COMPLEX_POLAR'(0.0, 0.0) if Z.MAG = 1.0 and
        --                                                Z.ARG = 0.0
        --         LOG(Z, BASE) = COMPLEX_POLAR'(1.0, 0.0) if Z.MAG = BASE and
        --                                                Z.ARG = 0.0
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        --         Z.MAG /= 0.0
        --         BASE > 0.0
        --         BASE /= 1.0
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        --         Error if Z.MAG = 0.0
        --         Error if BASE <= 0.0
        --         Error if BASE = 1.0
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function SIN (Z : in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns sine of Z
        -- Special values:
        --         SIN(MATH_CZERO) = MATH_CZERO
        --         SIN(Z) = MATH_CZERO if Z = COMPLEX'(MATH_PI, 0.0)
        -- Domain:
        --         Z in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         ABS(SIN(Z)) <= SQRT(SIN(Z.RE)*SIN(Z.RE) +
        --                                         SINH(Z.IM)*SINH(Z.IM))
        -- Notes:
        --         None

    function SIN (Z : in COMPLEX_POLAR ) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns principal value of sine of Z
        -- Special values:
        --         SIN(Z) = COMPLEX_POLAR'(0.0, 0.0) if Z.MAG = 0.0 and
        --                                            Z.ARG = 0.0
        --         SIN(Z) = COMPLEX_POLAR'(0.0, 0.0) if Z.MAG = MATH_PI and
        --                                            Z.ARG = 0.0
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function  COS (Z : in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns cosine of Z
        -- Special values:
        --         COS(Z) = MATH_CZERO if Z = COMPLEX'(MATH_PI_OVER_2, 0.0)
        --         COS(Z) = MATH_CZERO if Z = COMPLEX'(-MATH_PI_OVER_2, 0.0)
        -- Domain:
        --         Z in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         ABS(COS(Z)) <= SQRT(COS(Z.RE)*COS(Z.RE) +
        --                                         SINH(Z.IM)*SINH(Z.IM))
        -- Notes:
        --         None


    function  COS (Z : in COMPLEX_POLAR ) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns principal value of cosine of Z
        -- Special values:
        --         COS(Z) = COMPLEX_POLAR'(0.0, 0.0) if Z.MAG = MATH_PI_OVER_2
        --                                               and Z.ARG = 0.0
        --         COS(Z) = COMPLEX_POLAR'(0.0, 0.0) if Z.MAG = MATH_PI_OVER_2
        --                                               and Z.ARG = MATH_PI
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function SINH (Z : in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns hyperbolic sine of Z
        -- Special values:
        --         SINH(MATH_CZERO) = MATH_CZERO
        --         SINH(Z) = MATH_CZERO if Z.RE = 0.0 and Z.IM = MATH_PI
        --         SINH(Z) = MATH_CBASE_J if Z.RE = 0.0 and
        --                                               Z.IM = MATH_PI_OVER_2
        --         SINH(Z) = -MATH_CBASE_J if Z.RE = 0.0 and
        --                                               Z.IM = -MATH_PI_OVER_2
        -- Domain:
        --         Z in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         ABS(SINH(Z)) <= SQRT(SINH(Z.RE)*SINH(Z.RE) +
        --                                         SIN(Z.IM)*SIN(Z.IM))
        -- Notes:
        --         None

    function SINH (Z : in COMPLEX_POLAR ) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns principal value of hyperbolic sine of Z
        -- Special values:
        --         SINH(Z) = COMPLEX_POLAR'(0.0, 0.0) if Z.MAG = 0.0 and
        --                                            Z.ARG = 0.0
        --         SINH(Z) = COMPLEX_POLAR'(0.0, 0.0) if Z.MAG = MATH_PI and
        --                                            Z.ARG = MATH_PI_OVER_2
        --         SINH(Z) = COMPLEX_POLAR'(1.0, MATH_PI_OVER_2) if Z.MAG =
        --                         MATH_PI_OVER_2 and Z.ARG = MATH_PI_OVER_2
        --         SINH(Z) = COMPLEX_POLAR'(1.0, -MATH_PI_OVER_2) if Z.MAG =
        --                         MATH_PI_OVER_2 and Z.ARG = -MATH_PI_OVER_2
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function COSH (Z : in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns hyperbolic cosine of Z
        -- Special values:
        --         COSH(MATH_CZERO) = MATH_CBASE_1
        --         COSH(Z) = -MATH_CBASE_1 if Z.RE = 0.0 and Z.IM = MATH_PI
        --         COSH(Z) = MATH_CZERO if Z.RE = 0.0 and Z.IM = MATH_PI_OVER_2
        --         COSH(Z) = MATH_CZERO if Z.RE = 0.0 and Z.IM = -MATH_PI_OVER_2
        -- Domain:
        --         Z in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         ABS(COSH(Z)) <= SQRT(SINH(Z.RE)*SINH(Z.RE) +
        --                                         COS(Z.IM)*COS(Z.IM))
        -- Notes:
        --         None


    function COSH (Z : in COMPLEX_POLAR ) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns principal value of hyperbolic cosine of Z
        -- Special values:
        --         COSH(Z) = COMPLEX_POLAR'(1.0, 0.0) if Z.MAG = 0.0 and
        --                                            Z.ARG = 0.0
        --         COSH(Z) = COMPLEX_POLAR'(1.0, MATH_PI) if Z.MAG = MATH_PI and
        --                                            Z.ARG = MATH_PI_OVER_2
        --         COSH(Z) = COMPLEX_POLAR'(0.0, 0.0) if Z.MAG =
        --                        MATH_PI_OVER_2 and Z.ARG = MATH_PI_OVER_2
        --         COSH(Z) = COMPLEX_POLAR'(0.0, 0.0) if Z.MAG =
        --                        MATH_PI_OVER_2 and Z.ARG = -MATH_PI_OVER_2
        -- Domain:
        --         Z in COMPLEX_POLAR and Z.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if Z.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    --
    -- Arithmetic Operators
    --

    function "+" ( L: in COMPLEX;  R: in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns arithmetic addition of L and R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX
        --         R in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         "+"(Z) is mathematically unbounded
        -- Notes:
        --         None

    function "+" ( L: in REAL;     R: in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns arithmetic addition of L and R
        -- Special values:
        --         None
        -- Domain:
        --         L in REAL
        --         R in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         "+"(Z) is mathematically unbounded
        -- Notes:
        --         None

    function "+" ( L: in COMPLEX;  R: in REAL )    return COMPLEX;
        -- Purpose:
        --         Returns arithmetic addition of L and R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX
        --         R in REAL
        -- Error conditions:
        --         None
        -- Range:
        --         "+"(Z) is mathematically unbounded
        -- Notes:
        --         None

    function "+" ( L: in COMPLEX_POLAR; R: in COMPLEX_POLAR)
                                                        return COMPLEX_POLAR;
        -- Purpose:
        --         Returns arithmetic addition of L and R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX_POLAR and L.ARG /= -MATH_PI
        --         R in COMPLEX_POLAR and R.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if L.ARG = -MATH_PI
        --         Error if R.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None


    function "+" ( L: in REAL;  R: in COMPLEX_POLAR) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns arithmetic addition of L and R
        -- Special values:
        --         None
        -- Domain:
        --         L in REAL
        --         R in COMPLEX_POLAR and R.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if R.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function "+" ( L: in COMPLEX_POLAR;  R: in REAL) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns arithmetic addition of L and R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX_POLAR and L.ARG /= -MATH_PI
        --         R in REAL
        -- Error conditions:
        --         Error if L.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function "-" ( L: in COMPLEX;  R: in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns arithmetic subtraction of L minus R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX
        --         R in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         "-"(Z) is mathematically unbounded
        -- Notes:
        --         None

    function "-" ( L: in REAL;     R: in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns arithmetic subtraction of L minus R
        -- Special values:
        --         None
        -- Domain:
        --         L in REAL
        --         R in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         "-"(Z) is mathematically unbounded
        -- Notes:
        --         None

    function "-" ( L: in COMPLEX;  R: in REAL )    return COMPLEX;
        -- Purpose:
        --         Returns arithmetic subtraction of L minus R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX
        --         R in REAL
        -- Error conditions:
        --         None
        -- Range:
        --         "-"(Z) is mathematically unbounded
        -- Notes:
        --         None

    function "-" ( L: in COMPLEX_POLAR; R: in COMPLEX_POLAR)
                                                        return COMPLEX_POLAR;
        -- Purpose:
        --         Returns arithmetic subtraction of L minus R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX_POLAR and L.ARG /= -MATH_PI
        --         R in COMPLEX_POLAR and R.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if L.ARG = -MATH_PI
        --         Error if R.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function "-" ( L: in REAL;  R: in COMPLEX_POLAR) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns arithmetic subtraction of L minus R
        -- Special values:
        --         None
        -- Domain:
        --         L in REAL
        --         R in COMPLEX_POLAR and R.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if R.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None


    function "-" ( L: in COMPLEX_POLAR;  R: in REAL) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns arithmetic subtraction of L minus R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX_POLAR and L.ARG /= -MATH_PI
        --         R in REAL
        -- Error conditions:
        --         Error if L.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function "*" ( L: in COMPLEX;  R: in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns arithmetic multiplication of L and R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX
        --         R in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         "*"(Z) is mathematically unbounded
        -- Notes:
        --         None

    function "*" ( L: in REAL;  R: in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns arithmetic multiplication of L and R
        -- Special values:
        --         None
        -- Domain:
        --         L in REAL
        --         R in COMPLEX
        -- Error conditions:
        --         None
        -- Range:
        --         "*"(Z) is mathematically unbounded
        -- Notes:
        --         None

    function "*" ( L: in COMPLEX;  R: in REAL )  return COMPLEX;
        -- Purpose:
        --         Returns arithmetic multiplication of L and R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX
        --         R in REAL
        -- Error conditions:
        --         None

        -- Range:
        --         "*"(Z) is mathematically unbounded
        -- Notes:
        --         None

    function "*" ( L: in COMPLEX_POLAR; R: in COMPLEX_POLAR)
                                                        return COMPLEX_POLAR;
        -- Purpose:
        --         Returns arithmetic multiplication of L and R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX_POLAR and L.ARG /= -MATH_PI
        --         R in COMPLEX_POLAR and R.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if L.ARG = -MATH_PI
        --         Error if R.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function "*" ( L: in REAL;  R: in COMPLEX_POLAR) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns arithmetic multiplication of L and R
        -- Special values:
        --         None
        -- Domain:
        --         L in REAL
        --         R in COMPLEX_POLAR and R.ARG /= -MATH_PI
        -- Error conditions:
        --         Error if R.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function "*" ( L: in COMPLEX_POLAR;  R: in REAL) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns arithmetic multiplication of L and R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX_POLAR and L.ARG /= -MATH_PI
        --         R in REAL
        -- Error conditions:
        --         Error if L.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None


    function "/" ( L: in COMPLEX;  R: in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns arithmetic division of L by R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX
        --         R in COMPLEX and R /= MATH_CZERO
        -- Error conditions:
        --         Error if R = MATH_CZERO
        -- Range:
        --         "/"(Z) is mathematically unbounded
        -- Notes:
        --         None

    function "/" ( L: in REAL;  R: in COMPLEX ) return COMPLEX;
        -- Purpose:
        --         Returns arithmetic division of L by R
        -- Special values:
        --         None
        -- Domain:
        --         L in REAL
        --         R in COMPLEX and R /= MATH_CZERO
        -- Error conditions:
        --         Error if R = MATH_CZERO
        -- Range:
        --         "/"(Z) is mathematically unbounded
        -- Notes:
        --         None

    function "/" ( L: in COMPLEX;  R: in REAL )    return COMPLEX;
        -- Purpose:
        --         Returns arithmetic division of L by R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX
        --         R in REAL and R /= 0.0
        -- Error conditions:
        --         Error if R = 0.0
        -- Range:
        --         "/"(Z) is mathematically unbounded
        -- Notes:
        --         None

    function "/" ( L: in COMPLEX_POLAR; R: in COMPLEX_POLAR)
                                                        return COMPLEX_POLAR;
        -- Purpose:
        --         Returns arithmetic division of L by R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX_POLAR and L.ARG /= -MATH_PI
        --         R in COMPLEX_POLAR and R.ARG /= -MATH_PI
        --         R.MAG > 0.0
        -- Error conditions:
        --         Error if R.MAG <= 0.0
        --         Error if L.ARG = -MATH_PI
        --         Error if R.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function "/" ( L: in REAL;  R: in COMPLEX_POLAR) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns arithmetic division of L by R
        -- Special values:
        --         None
        -- Domain:
        --         L in REAL
        --         R in COMPLEX_POLAR and R.ARG /= -MATH_PI
        --         R.MAG > 0.0
        -- Error conditions:
        --         Error if R.MAG <= 0.0
        --         Error if R.ARG = -MATH_PI
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None

    function "/" ( L: in COMPLEX_POLAR;  R: in REAL) return COMPLEX_POLAR;
        -- Purpose:
        --         Returns arithmetic division of L by R
        -- Special values:
        --         None
        -- Domain:
        --         L in COMPLEX_POLAR and L.ARG /= -MATH_PI
        --         R /= 0.0
        -- Error conditions:
        --         Error if L.ARG = -MATH_PI
        --         Error if R = 0.0
        -- Range:
        --         result.MAG >= 0.0
        --         -MATH_PI < result.ARG <= MATH_PI
        -- Notes:
        --         None
end  MATH_COMPLEX;




------------------------------------------------------------------------
--
-- Copyright 1996 by IEEE. All rights reserved.
--
-- This source file is an informative part of IEEE Std 1076.2-1996, IEEE Standard 
-- VHDL Mathematical Packages. This source file may not be copied, sold, or 
-- included with software that is sold without written permission from the IEEE
-- Standards Department. This source file may be used to implement this standard 
-- and may be distributed in compiled form in any manner so long as the 
-- compiled form does not allow direct decompilation of the original source file.
-- This source file may be copied for individual use between licensed users. 
-- This source file is provided on an AS IS basis. The IEEE disclaims ANY 
-- WARRANTY EXPRESS OR IMPLIED INCLUDING ANY WARRANTY OF MERCHANTABILITY 
-- AND FITNESS FOR USE FOR A PARTICULAR PURPOSE. The user of the source 
-- file shall indemnify and hold IEEE harmless from any damages or liability 
-- arising out of the use thereof.
--
-- Title:       Standard VHDL Mathematical Packages (IEEE Std 1076.2-1996,
--              MATH_COMPLEX)
--
-- Library:     This package shall be compiled into a library
--              symbolically named IEEE.
--
-- Developers:  IEEE DASC VHDL Mathematical Packages Working Group
--
-- Purpose:     This package body is a nonnormative implementation of the 
--              functionality defined in the MATH_COMPLEX package declaration.
--
-- Limitation:  The values generated by the functions in this package may
--              vary from platform to platform, and the precision of results
--              is only guaranteed to be the minimum required by IEEE Std 1076
--              -1993.
--
-- Notes:
--              The "package declaration" defines the types, subtypes, and
--              declarations of MATH_COMPLEX.
--              The standard mathematical definition and conventional meaning
--              of the mathematical functions that are part of this standard
--              represent the formal semantics of the implementation of the
--              MATH_COMPLEX package declaration.  The purpose of the
--              MATH_COMPLEX package body is to clarify such semantics and
--              provide a guideline for implementations to verify their
--              implementation of MATH_COMPLEX.  Tool developers may choose to
--              implement the package body in the most efficient manner
--              available to them.
--
-- -----------------------------------------------------------------------------
-- Version    : 1.5
-- Date       : 24 July 1996
-- -----------------------------------------------------------------------------
library IEEE;
use IEEE.MATH_REAL.all;

package body MATH_COMPLEX is

    --
    -- Equality and Inequality Operators for COMPLEX_POLAR
    --
    function "=" ( L: in COMPLEX_POLAR;  R: in COMPLEX_POLAR ) return BOOLEAN
                                                                         is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns FALSE on error
    begin
        -- Check validity of input arguments
        if ( L.ARG = -MATH_PI ) then
                assert FALSE
                            report "L.ARG = -MATH_PI in =(L,R)"
                            severity ERROR;
                return FALSE;
        end if;

        if ( R.ARG = -MATH_PI ) then
                assert FALSE
                            report "R.ARG = -MATH_PI in =(L,R)"
                            severity ERROR;
                return FALSE;
        end if;

        -- Get special values
        if ( L.MAG = 0.0 and R.MAG = 0.0 ) then
                return TRUE;
        end if;

        -- Get value for general case
        if ( L.MAG = R.MAG and L.ARG = R.ARG ) then
                return TRUE;
        end if;

        return FALSE;
    end "=";


    function "/=" ( L: in COMPLEX_POLAR;  R: in COMPLEX_POLAR ) return BOOLEAN
                                                                         is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns FALSE on error
    begin
        -- Check validity of input arguments
        if ( L.ARG = -MATH_PI ) then
                assert FALSE
                            report "L.ARG = -MATH_PI in /=(L,R)"
                            severity ERROR;
                return FALSE;
        end if;

        if ( R.ARG = -MATH_PI ) then
                assert FALSE
                            report "R.ARG = -MATH_PI in /=(L,R)"
                            severity ERROR;
                return FALSE;
        end if;

        -- Get special values
        if ( L.MAG = 0.0 and R.MAG = 0.0 ) then
                return FALSE;
        end if;

        -- Get value for general case
        if ( L.MAG = R.MAG and L.ARG = R.ARG ) then
                return FALSE;
        end if;

        return TRUE;
    end "/=";

    --
    -- Other Functions Start Here
    --

    function CMPLX(X: in REAL;  Y: in REAL := 0.0 ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
    begin
        return COMPLEX'(X, Y);
    end CMPLX;


    function GET_PRINCIPAL_VALUE(X: in REAL ) return PRINCIPAL_VALUE is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
        variable TEMP: REAL;
    begin
        -- Check if already a principal value
        if ( X > -MATH_PI and X <= MATH_PI ) then
                return PRINCIPAL_VALUE'(X);
        end if;

        -- Get principal value
        TEMP := X;
        while ( TEMP <= -MATH_PI ) loop
                TEMP := TEMP + MATH_2_PI;
        end loop;
        while (TEMP > MATH_PI ) loop
                TEMP := TEMP - MATH_2_PI;
        end loop;

        return PRINCIPAL_VALUE'(TEMP);
    end GET_PRINCIPAL_VALUE;

    function COMPLEX_TO_POLAR(Z: in COMPLEX ) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
        variable TEMP: REAL;
    begin
        -- Get value for special cases
        if ( Z.RE = 0.0 ) then
            if ( Z.IM = 0.0 ) then
                return COMPLEX_POLAR'(0.0, 0.0);
            elsif ( Z.IM > 0.0 ) then
                return COMPLEX_POLAR'(Z.IM, MATH_PI_OVER_2);
            else
                return COMPLEX_POLAR'(-Z.IM, -MATH_PI_OVER_2);
            end if;
        end if;

        if ( Z.IM = 0.0 ) then
            if ( Z.RE = 0.0 ) then
                return COMPLEX_POLAR'(0.0, 0.0);
            elsif ( Z.RE > 0.0 ) then
                return COMPLEX_POLAR'(Z.RE, 0.0);
            else
                return COMPLEX_POLAR'(-Z.RE, MATH_PI);
            end if;
        end if;

        -- Get principal value for general case
        TEMP := ARCTAN(Z.IM, Z.RE);

        return COMPLEX_POLAR'(SQRT(Z.RE*Z.RE + Z.IM*Z.IM),
                                                 GET_PRINCIPAL_VALUE(TEMP));
    end COMPLEX_TO_POLAR;

    function POLAR_TO_COMPLEX(Z: in COMPLEX_POLAR ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns MATH_CZERO on error
    begin
        -- Check validity of input arguments
        if ( Z.ARG = -MATH_PI ) then
                assert FALSE
                       report "Z.ARG = -MATH_PI in POLAR_TO_COMPLEX(Z)"
                       severity ERROR;
                return MATH_CZERO;
        end if;

        -- Get value for general case
        return COMPLEX'( Z.MAG*COS(Z.ARG), Z.MAG*SIN(Z.ARG) );
    end POLAR_TO_COMPLEX;


    function "ABS"(Z: in COMPLEX ) return POSITIVE_REAL is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) ABS(Z) = SQRT(Z.RE*Z.RE + Z.IM*Z.IM)

    begin
        -- Get value for general case
        return POSITIVE_REAL'(SQRT(Z.RE*Z.RE + Z.IM*Z.IM));
    end "ABS";

    function "ABS"(Z: in COMPLEX_POLAR ) return POSITIVE_REAL is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) ABS(Z) = Z.MAG
        --        b) Returns 0.0 on error

    begin
        -- Check validity of input arguments
        if ( Z.ARG = -MATH_PI ) then
                  assert FALSE
                            report "Z.ARG = -MATH_PI in ABS(Z)"
                            severity ERROR;
                  return 0.0;
        end if;

        -- Get value for general case
        return Z.MAG;
    end "ABS";


    function ARG(Z: in COMPLEX ) return PRINCIPAL_VALUE is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) ARG(Z) = ARCTAN(Z.IM, Z.RE)

        variable ZTEMP : COMPLEX_POLAR;
    begin
        -- Get value for general case
        ZTEMP := COMPLEX_TO_POLAR(Z);
        return ZTEMP.ARG;
    end ARG;

    function ARG(Z: in COMPLEX_POLAR ) return PRINCIPAL_VALUE is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) ARG(Z) = Z.ARG
        --        b) Returns 0.0 on error

    begin
        -- Check validity of input arguments
        if ( Z.ARG = -MATH_PI ) then
                  assert FALSE
                            report "Z.ARG = -MATH_PI in ARG(Z)"
                            severity ERROR;
                  return 0.0;
        end if;

        -- Get value for general case
        return Z.ARG;
    end ARG;

    function "-" (Z: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns -x -jy for Z = x + jy
    begin
        -- Get value for general case
        return COMPLEX'(-Z.RE, -Z.IM);
    end "-";

    function "-" (Z: in COMPLEX_POLAR ) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns (Z.MAG, Z.ARG + MATH_PI)
        --        b) Returns Z on error
        variable TEMP: REAL;
    begin
        -- Check validity of input arguments
        if ( Z.ARG = -MATH_PI ) then
                  assert FALSE
                            report "Z.ARG = -MATH_PI in -(Z)"
                            severity ERROR;
                  return Z;
        end if;

        -- Get principal value for general case
        TEMP := REAL'(Z.ARG) + MATH_PI;

        return COMPLEX_POLAR'(Z.MAG, GET_PRINCIPAL_VALUE(TEMP));
    end "-";

    function CONJ (Z: in COMPLEX) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns x - jy for Z = x + jy
    begin
        -- Get value for general case
        return COMPLEX'(Z.RE, -Z.IM);
    end CONJ;

    function CONJ (Z: in COMPLEX_POLAR) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX conjugate (Z.MAG, -Z.ARG)
        --        b) Returns Z on error
        --
        variable TEMP: PRINCIPAL_VALUE;
    begin
        -- Check validity of input arguments
        if ( Z.ARG = -MATH_PI ) then
                  assert FALSE
                            report "Z.ARG = -MATH_PI in CONJ(Z)"
                            severity ERROR;
                  return Z;
        end if;

        -- Get principal value for general case
        if ( Z.ARG = MATH_PI or Z.ARG = 0.0 ) then
                TEMP := Z.ARG;
        else
                TEMP := -Z.ARG;
        end if;

         return COMPLEX_POLAR'(Z.MAG, TEMP);
    end CONJ;

    function SQRT(Z: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
        variable ZTEMP : COMPLEX_POLAR;
        variable ZOUT : COMPLEX;
        variable TMAG : REAL;
        variable TARG : REAL;
    begin
        -- Get value for special cases
        if ( Z = MATH_CZERO ) then
                return MATH_CZERO;
        end if;

        -- Get value for general case
        ZTEMP := COMPLEX_TO_POLAR(Z);
        TMAG := SQRT(ZTEMP.MAG);
        TARG := 0.5*ZTEMP.ARG;

        if ( COS(TARG) > 0.0 ) then
                ZOUT.RE := TMAG*COS(TARG);
                ZOUT.IM := TMAG*SIN(TARG);
                return ZOUT;
        end if;

        if ( COS(TARG) < 0.0 ) then
                ZOUT.RE := TMAG*COS(TARG + MATH_PI);
                ZOUT.IM := TMAG*SIN(TARG + MATH_PI);
                return ZOUT;
        end if;

        if ( SIN(TARG) > 0.0 ) then
                ZOUT.RE := 0.0;
                ZOUT.IM := TMAG*SIN(TARG);
                return ZOUT;
        end if;

        ZOUT.RE := 0.0;
        ZOUT.IM := TMAG*SIN(TARG + MATH_PI);
        return ZOUT;
    end SQRT;

    function SQRT(Z: in COMPLEX_POLAR ) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns Z on error

        variable ZOUT : COMPLEX_POLAR;
        variable TMAG : REAL;
        variable TARG : REAL;
    begin
        -- Check validity of input arguments
        if ( Z.ARG = -MATH_PI ) then
                  assert FALSE
                            report "Z.ARG = -MATH_PI in SQRT(Z)"
                            severity ERROR;
                  return Z;
        end if;

        -- Get value for special cases
        if ( Z.MAG = 0.0 and Z.ARG = 0.0 ) then
                return Z;
        end if;

        -- Get principal value for general case
        TMAG := SQRT(Z.MAG);
        TARG := 0.5*Z.ARG;

        ZOUT.MAG := POSITIVE_REAL'(TMAG);

        if ( COS(TARG) < 0.0 ) then
                TARG := TARG + MATH_PI;
        end if;

        if ( (COS(TARG) = 0.0) and (SIN(TARG) < 0.0) ) then
                TARG := TARG + MATH_PI;
        end if;

        ZOUT.ARG := GET_PRINCIPAL_VALUE(TARG);
        return ZOUT;
    end SQRT;

    function EXP(Z: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None

        variable TEMP: REAL;
    begin
        -- Get value for special cases
        if ( Z = MATH_CZERO ) then
                return MATH_CBASE_1;
        end if;

        if ( Z.RE = 0.0 ) then
                if ( Z.IM = MATH_PI or Z.IM = -MATH_PI ) then
                        return COMPLEX'(-1.0, 0.0);
                end if;

                if ( Z.IM = MATH_PI_OVER_2 ) then
                        return MATH_CBASE_J;
                end if;

                if ( Z.IM = -MATH_PI_OVER_2 ) then
                        return COMPLEX'(0.0, -1.0);
                end if;
        end if;

        -- Get value for general case
        TEMP := EXP(Z.RE);
        return COMPLEX'(TEMP*COS(Z.IM), TEMP*SIN(Z.IM));
    end EXP;

    function EXP(Z: in COMPLEX_POLAR ) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns Z on error

        variable ZTEMP : COMPLEX;
        variable temp: REAL;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( Z.ARG = -MATH_PI ) then
                  assert FALSE
                            report "Z.ARG = -MATH_PI in EXP(Z)"
                            severity ERROR;
                  return Z;
        end if;

        -- Get value for special cases
        if ( Z.MAG = 0.0 and Z.ARG = 0.0 ) then
                return COMPLEX_POLAR'(1.0, 0.0);
        end if;

        if ( Z.MAG = MATH_PI and (Z.ARG = MATH_PI_OVER_2 or
                                                 Z.ARG = -MATH_PI_OVER_2 )) then
                return COMPLEX_POLAR'(1.0, MATH_PI);
        end if;

        if ( Z.MAG = MATH_PI_OVER_2 ) then
                if ( Z.ARG = MATH_PI_OVER_2 ) then
                        return COMPLEX_POLAR'(1.0, MATH_PI_OVER_2);
                end if;

                if ( Z.ARG = -MATH_PI_OVER_2 ) then
                        return COMPLEX_POLAR'(1.0, -MATH_PI_OVER_2);
                end if;
        end if;

        -- Get principal value for general case
        ZTEMP := POLAR_TO_COMPLEX(Z);
        ZOUT.MAG := POSITIVE_REAL'(EXP(ZTEMP.RE));
        ZOUT.ARG := GET_PRINCIPAL_VALUE(ZTEMP.IM);

        return ZOUT;
    end EXP;

    function LOG(Z: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX'(REAL'LOW, 0.0) on error

        variable ZTEMP : COMPLEX_POLAR;
        variable TEMP : REAL;
    begin
        -- Check validity of input arguments
        if ( Z.RE = 0.0  and Z.IM = 0.0 ) then
                assert FALSE
                        report "Z.RE = 0.0 and Z.IM = 0.0 in LOG(Z)"
                        severity ERROR;
                return COMPLEX'(REAL'LOW, 0.0);
        end if;

        -- Get value for special cases
        if ( Z.IM = 0.0 ) then
                if ( Z.RE = -1.0 ) then
                        return COMPLEX'(0.0, MATH_PI);
                end if;
                if ( Z.RE = MATH_E ) then
                        return MATH_CBASE_1;
                end if;
                if ( Z.RE = 1.0 ) then
                        return MATH_CZERO;
                end if;
        end if;

        if ( Z.RE = 0.0 ) then
                if (Z.IM = 1.0) then
                        return COMPLEX'(0.0, MATH_PI_OVER_2);
                end if;
                if (Z.IM = -1.0) then
                        return COMPLEX'(0.0, -MATH_PI_OVER_2);
                end if;
        end if;

        -- Get value for general case
        ZTEMP := COMPLEX_TO_POLAR(Z);
        TEMP := LOG(ZTEMP.MAG);
        return COMPLEX'(TEMP, ZTEMP.ARG);
    end LOG;

    function LOG2(Z: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX'(REAL'LOW, 0.0) on error

        variable ZTEMP : COMPLEX_POLAR;
        variable TEMP : REAL;
    begin

        -- Check validity of input arguments
        if ( Z.RE = 0.0  and Z.IM = 0.0 ) then
                assert FALSE
                        report "Z.RE = 0.0 and Z.IM = 0.0 in LOG2(Z)"
                        severity ERROR;
                return COMPLEX'(REAL'LOW, 0.0);
        end if;

        -- Get value for special cases
        if ( Z.IM = 0.0 ) then
                if ( Z.RE = 2.0 ) then
                        return MATH_CBASE_1;
                end if;
                if ( Z.RE = 1.0 ) then
                        return MATH_CZERO;
                end if;
        end if;

        -- Get value for general case
        ZTEMP := COMPLEX_TO_POLAR(Z);
        TEMP := MATH_LOG2_OF_E*LOG(ZTEMP.MAG);
        return COMPLEX'(TEMP, MATH_LOG2_OF_E*ZTEMP.ARG);
    end LOG2;

    function LOG10(Z: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX'(REAL'LOW, 0.0) on error

        variable ZTEMP : COMPLEX_POLAR;
        variable TEMP : REAL;
    begin
        -- Check validity of input arguments
        if ( Z.RE = 0.0  and Z.IM = 0.0 ) then
                assert FALSE
                        report "Z.RE = 0.0 and Z.IM = 0.0 in LOG10(Z)"
                        severity ERROR;
                return COMPLEX'(REAL'LOW, 0.0);
        end if;

        -- Get value for special cases
        if ( Z.IM = 0.0 ) then
                if ( Z.RE = 10.0 ) then
                        return MATH_CBASE_1;
                end if;
                if ( Z.RE = 1.0 ) then
                        return MATH_CZERO;
                end if;
        end if;

        -- Get value for general case
        ZTEMP := COMPLEX_TO_POLAR(Z);
        TEMP := MATH_LOG10_OF_E*LOG(ZTEMP.MAG);
        return COMPLEX'(TEMP, MATH_LOG10_OF_E*ZTEMP.ARG);
    end LOG10;


    function LOG(Z: in COMPLEX_POLAR ) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR(REAL'HIGH, MATH_PI) on error

        variable ZTEMP : COMPLEX;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( Z.MAG <= 0.0 ) then
                assert FALSE
                        report "Z.MAG <= 0.0 in LOG(Z)"
                        severity ERROR;
                return COMPLEX_POLAR'(REAL'HIGH, MATH_PI);
        end if;

        if ( Z.ARG = -MATH_PI ) then
                  assert FALSE
                            report "Z.ARG = -MATH_PI in LOG(Z)"
                            severity ERROR;
                return COMPLEX_POLAR'(REAL'HIGH, MATH_PI);
        end if;

        -- Compute value for special cases
        if (Z.MAG = 1.0 ) then
                if ( Z.ARG = 0.0 ) then
                        return COMPLEX_POLAR'(0.0, 0.0);
                end if;

                if ( Z.ARG = MATH_PI ) then
                        return COMPLEX_POLAR'(MATH_PI, MATH_PI_OVER_2);
                end if;

                if ( Z.ARG = MATH_PI_OVER_2 ) then
                        return COMPLEX_POLAR'(MATH_PI_OVER_2, MATH_PI_OVER_2);
                end if;

                if ( Z.ARG = -MATH_PI_OVER_2 ) then
                        return COMPLEX_POLAR'(MATH_PI_OVER_2, -MATH_PI_OVER_2);
                end if;
        end if;

        if ( Z.MAG = MATH_E and Z.ARG = 0.0 ) then
                return COMPLEX_POLAR'(1.0, 0.0);
        end if;

        -- Compute value for general case
        ZTEMP.RE := LOG(Z.MAG);
        ZTEMP.IM := Z.ARG;
        ZOUT := COMPLEX_TO_POLAR(ZTEMP);
        return ZOUT;
    end LOG;



    function LOG2(Z: in COMPLEX_POLAR ) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR(REAL'HIGH, MATH_PI) on error

        variable ZTEMP : COMPLEX;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( Z.MAG <= 0.0 ) then
                assert FALSE
                        report "Z.MAG <= 0.0 in LOG2(Z)"
                        severity ERROR;
                return COMPLEX_POLAR'(REAL'HIGH, MATH_PI);
        end if;

        if ( Z.ARG = -MATH_PI ) then
                  assert FALSE
                            report "Z.ARG = -MATH_PI in LOG2(Z)"
                            severity ERROR;
                return COMPLEX_POLAR'(REAL'HIGH, MATH_PI);
        end if;

        -- Compute value for special cases
        if (Z.MAG = 1.0 and Z.ARG = 0.0 ) then
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        if ( Z.MAG = 2.0 and Z.ARG = 0.0 ) then
                return COMPLEX_POLAR'(1.0, 0.0);
        end if;

        -- Compute value for general case
        ZTEMP.RE := MATH_LOG2_OF_E*LOG(Z.MAG);
        ZTEMP.IM := MATH_LOG2_OF_E*Z.ARG;
        ZOUT := COMPLEX_TO_POLAR(ZTEMP);
        return ZOUT;
    end LOG2;

    function LOG10(Z: in COMPLEX_POLAR ) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR(REAL'HIGH, MATH_PI) on error
        variable ZTEMP : COMPLEX;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( Z.MAG <= 0.0 ) then
                assert FALSE
                        report "Z.MAG <= 0.0 in LOG10(Z)"
                        severity ERROR;
                return COMPLEX_POLAR'(REAL'HIGH, MATH_PI);
        end if;


        if ( Z.ARG = -MATH_PI ) then
                  assert FALSE
                           report "Z.ARG = -MATH_PI in LOG10(Z)"
                           severity ERROR;
                return COMPLEX_POLAR'(REAL'HIGH, MATH_PI);
        end if;

        -- Compute value for special cases
        if (Z.MAG = 1.0 and Z.ARG = 0.0 ) then
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        if ( Z.MAG = 10.0 and Z.ARG = 0.0 ) then
                return COMPLEX_POLAR'(1.0, 0.0);
        end if;

        -- Compute value for general case
        ZTEMP.RE := MATH_LOG10_OF_E*LOG(Z.MAG);
        ZTEMP.IM := MATH_LOG10_OF_E*Z.ARG;
        ZOUT := COMPLEX_TO_POLAR(ZTEMP);
        return ZOUT;
    end LOG10;

    function LOG(Z: in COMPLEX; BASE: in REAL ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX'(REAL'LOW, 0.0) on error

        variable ZTEMP : COMPLEX_POLAR;
        variable TEMPRE : REAL;
        variable TEMPIM : REAL;
    begin
        -- Check validity of input arguments
        if ( Z.RE = 0.0  and Z.IM = 0.0 ) then
                assert FALSE
                        report "Z.RE = 0.0 and Z.IM = 0.0 in LOG(Z,BASE)"
                        severity ERROR;
                return COMPLEX'(REAL'LOW, 0.0);
        end if;

        if ( BASE <= 0.0 or BASE = 1.0 ) then
                assert FALSE
                        report "BASE <= 0.0 or BASE = 1.0 in LOG(Z,BASE)"
                        severity ERROR;
                return COMPLEX'(REAL'LOW, 0.0);
        end if;

        -- Get value for special cases
        if ( Z.IM = 0.0 ) then
                if ( Z.RE = BASE ) then
                        return MATH_CBASE_1;
                end if;
                if ( Z.RE = 1.0 ) then
                        return MATH_CZERO;
                end if;
        end if;

        -- Get value for general case
        ZTEMP := COMPLEX_TO_POLAR(Z);
        TEMPRE := LOG(ZTEMP.MAG, BASE);
        TEMPIM := ZTEMP.ARG/LOG(BASE);
        return COMPLEX'(TEMPRE, TEMPIM);
    end LOG;

    function LOG(Z: in COMPLEX_POLAR; BASE: in REAL ) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR(REAL'HIGH, MATH_PI) on error

        variable ZTEMP : COMPLEX;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( Z.MAG <= 0.0 ) then
                assert FALSE
                        report "Z.MAG <= 0.0 in LOG(Z,BASE)"
                        severity ERROR;
                return COMPLEX_POLAR'(REAL'HIGH, MATH_PI);
        end if;

        if ( BASE <= 0.0 or BASE = 1.0 ) then
                assert FALSE
                        report "BASE <= 0.0 or BASE = 1.0 in LOG(Z,BASE)"
                        severity ERROR;
                return COMPLEX_POLAR'(REAL'HIGH, MATH_PI);
        end if;

        if ( Z.ARG = -MATH_PI ) then
                assert FALSE
                           report "Z.ARG = -MATH_PI in LOG(Z,BASE)"
                           severity ERROR;
                return COMPLEX_POLAR'(REAL'HIGH, MATH_PI);
        end if;

        -- Compute value for special cases
        if (Z.MAG = 1.0 and Z.ARG = 0.0 ) then
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        if ( Z.MAG = BASE and Z.ARG = 0.0 ) then
                return COMPLEX_POLAR'(1.0, 0.0);
        end if;

        -- Compute value for general case
        ZTEMP.RE := LOG(Z.MAG, BASE);
        ZTEMP.IM := Z.ARG/LOG(BASE);
        ZOUT := COMPLEX_TO_POLAR(ZTEMP);
        return ZOUT;
    end LOG;


    function SIN(Z: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
    begin
        -- Get value for special cases
        if ( Z.IM = 0.0 ) then
                if ( Z.RE = 0.0 or Z.RE = MATH_PI) then
                        return MATH_CZERO;
                end if;
        end if;

        -- Get value for general case
        return COMPLEX'(SIN(Z.RE)*COSH(Z.IM), COS(Z.RE)*SINH(Z.IM));
    end SIN;

    function SIN(Z: in COMPLEX_POLAR ) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR(0.0, 0.0) on error

        variable Z1, Z2 : COMPLEX;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( Z.ARG = -MATH_PI ) then
                assert FALSE
                            report "Z.ARG = -MATH_PI in SIN(Z)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Compute value for special cases
        if ( Z.MAG = 0.0 and Z.ARG = 0.0 ) then
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        if ( Z.MAG = MATH_PI and Z.ARG = 0.0 ) then
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Compute value for general case
        Z1 := POLAR_TO_COMPLEX(Z);
        Z2 := COMPLEX'(SIN(Z1.RE)*COSH(Z1.IM), COS(Z1.RE)*SINH(Z1.IM));
        ZOUT := COMPLEX_TO_POLAR(Z2);
        return ZOUT;
    end SIN;

    function COS(Z: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
    begin


        -- Get value for special cases
        if ( Z.IM = 0.0 ) then
                if ( Z.RE = MATH_PI_OVER_2 or Z.RE = -MATH_PI_OVER_2) then
                        return MATH_CZERO;
                end if;
        end if;

        -- Get value for general case
        return COMPLEX'(COS(Z.RE)*COSH(Z.IM), -SIN(Z.RE)*SINH(Z.IM));
    end COS;

    function COS(Z: in COMPLEX_POLAR ) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR(0.0, 0.0) on error

        variable Z1, Z2 : COMPLEX;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( Z.ARG = -MATH_PI ) then
                assert FALSE
                            report "Z.ARG = -MATH_PI in COS(Z)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Compute value for special cases
        if ( Z.MAG = MATH_PI_OVER_2 and Z.ARG = 0.0 ) then
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        if ( Z.MAG = MATH_PI_OVER_2 and Z.ARG = MATH_PI ) then
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Compute value for general case
        Z1 := POLAR_TO_COMPLEX(Z);
        Z2 := COMPLEX'(COS(Z1.RE)*COSH(Z1.IM), -SIN(Z1.RE)*SINH(Z1.IM));
        ZOUT := COMPLEX_TO_POLAR(Z2);
        return ZOUT;
    end COS;

    function SINH(Z: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
    begin
        -- Get value for special cases
        if ( Z.RE = 0.0 ) then
                if ( Z.IM = 0.0 or Z.IM = MATH_PI ) then
                        return MATH_CZERO;
                end if;



                if ( Z.IM = MATH_PI_OVER_2 ) then
                        return MATH_CBASE_J;
                end if;

                if ( Z.IM = -MATH_PI_OVER_2 ) then
                        return -MATH_CBASE_J;
                end if;
        end if;

        -- Get value for general case
        return COMPLEX'(SINH(Z.RE)*COS(Z.IM), COSH(Z.RE)*SIN(Z.IM));
    end SINH;

    function SINH(Z: in COMPLEX_POLAR ) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR(0.0, 0.0) on error

        variable Z1, Z2 : COMPLEX;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( Z.ARG = -MATH_PI ) then
                assert FALSE
                            report "Z.ARG = -MATH_PI in SINH(Z)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Compute value for special cases
        if ( Z.MAG = 0.0 and Z.ARG = 0.0 ) then
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        if ( Z.MAG = MATH_PI and Z.ARG = MATH_PI_OVER_2 ) then
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        if ( Z.MAG = MATH_PI_OVER_2 and Z.ARG = MATH_PI_OVER_2 ) then
                return COMPLEX_POLAR'(1.0, MATH_PI_OVER_2);
        end if;

        if ( Z.MAG = MATH_PI_OVER_2 and Z.ARG = -MATH_PI_OVER_2 ) then
                return COMPLEX_POLAR'(1.0, -MATH_PI_OVER_2);
        end if;

        -- Compute value for general case
        Z1 := POLAR_TO_COMPLEX(Z);
        Z2 := COMPLEX'(SINH(Z1.RE)*COS(Z1.IM), COSH(Z1.RE)*SIN(Z1.IM));
        ZOUT := COMPLEX_TO_POLAR(Z2);
        return ZOUT;
    end SINH;


    function COSH(Z: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
    begin
        -- Get value for special cases
        if ( Z.RE = 0.0 ) then
                if ( Z.IM = 0.0 ) then
                        return MATH_CBASE_1;
                end if;

                if ( Z.IM = MATH_PI ) then
                        return -MATH_CBASE_1;
                end if;

                if ( Z.IM = MATH_PI_OVER_2 or Z.IM = -MATH_PI_OVER_2 ) then
                        return MATH_CZERO;
                end if;
        end if;

        -- Get value for general case
        return COMPLEX'(COSH(Z.RE)*COS(Z.IM), SINH(Z.RE)*SIN(Z.IM));
    end COSH;

    function COSH(Z: in COMPLEX_POLAR ) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR(0.0, 0.0) on error

        variable Z1, Z2 : COMPLEX;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( Z.ARG = -MATH_PI ) then
                assert FALSE
                            report "Z.ARG = -MATH_PI in COSH(Z)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Compute value for special cases
        if ( Z.MAG = 0.0 and Z.ARG = 0.0 ) then
                return COMPLEX_POLAR'(1.0, 0.0);
        end if;

        if ( Z.MAG = MATH_PI and Z.ARG = MATH_PI_OVER_2 ) then
                return COMPLEX_POLAR'(1.0, MATH_PI);
        end if;

        if ( Z.MAG = MATH_PI_OVER_2 and Z.ARG = MATH_PI_OVER_2 ) then
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        if ( Z.MAG = MATH_PI_OVER_2 and Z.ARG = -MATH_PI_OVER_2 ) then
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Compute value for general case
        Z1 := POLAR_TO_COMPLEX(Z);
        Z2 := COMPLEX'(COSH(Z1.RE)*COS(Z1.IM), SINH(Z1.RE)*SIN(Z1.IM));
        ZOUT := COMPLEX_TO_POLAR(Z2);
        return ZOUT;
    end COSH;


    --
    -- Arithmetic Operators
    --
    function "+" ( L: in COMPLEX;  R: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
    begin
        return COMPLEX'(L.RE + R.RE, L.IM + R.IM);
    end "+";

    function "+" ( L: in REAL; R: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
    begin
        return COMPLEX'(L + R.RE, R.IM);
    end "+";

    function "+" ( L: in COMPLEX;  R: in REAL )    return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
    begin
        return COMPLEX'(L.RE + R, L.IM);
    end "+";

    function "+" (L: in COMPLEX_POLAR; R: in COMPLEX_POLAR)
                                                        return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR'(0.0, 0.0) on error
        --
        variable ZL, ZR : COMPLEX;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( L.ARG = -MATH_PI ) then
                assert FALSE
                            report "L.ARG = -MATH_PI in +(L,R)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;


        if ( R.ARG = -MATH_PI ) then
                assert FALSE
                            report "R.ARG = -MATH_PI in +(L,R)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Get principal value
        ZL := POLAR_TO_COMPLEX( L );
        ZR := POLAR_TO_COMPLEX( R );
        ZOUT := COMPLEX_TO_POLAR(COMPLEX'(ZL.RE + ZR.RE, ZL.IM +ZR.IM));
        return ZOUT;
    end "+";

    function "+" ( L: in REAL;  R: in COMPLEX_POLAR) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR'(0.0, 0.0) on error
        variable ZR : COMPLEX;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( R.ARG = -MATH_PI ) then
                assert FALSE
                            report "R.ARG = -MATH_PI in +(L,R)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Get principal value
        ZR := POLAR_TO_COMPLEX( R );
        ZOUT := COMPLEX_TO_POLAR(COMPLEX'(L + ZR.RE, ZR.IM));
        return ZOUT;
    end "+";

    function "+" ( L: in COMPLEX_POLAR;  R: in REAL) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR'(0.0, 0.0) on error
        --
        variable ZL : COMPLEX;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( L.ARG = -MATH_PI ) then
                assert FALSE
                            report "L.ARG = -MATH_PI in +(L,R)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Get principal value
        ZL := POLAR_TO_COMPLEX( L );
        ZOUT := COMPLEX_TO_POLAR(COMPLEX'(ZL.RE + R, ZL.IM));
        return ZOUT;
    end "+";

    function "-" ( L: in COMPLEX;  R: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
    begin
        return COMPLEX'(L.RE - R.RE, L.IM - R.IM);
    end "-";

    function "-" ( L: in REAL;     R: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
    begin
        return COMPLEX'(L - R.RE, -1.0 * R.IM);
    end "-";

    function "-" ( L: in COMPLEX;  R: in REAL )    return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
    begin
        return COMPLEX'(L.RE - R, L.IM);
    end "-";

    function "-" ( L: in COMPLEX_POLAR; R: in COMPLEX_POLAR)
                                                        return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR'(0.0, 0.0) on error
        --
        variable ZL, ZR : COMPLEX;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( L.ARG = -MATH_PI ) then
                assert FALSE
                            report "L.ARG = -MATH_PI in -(L,R)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        if ( R.ARG = -MATH_PI ) then
                assert FALSE
                            report "R.ARG = -MATH_PI in -(L,R)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;
        -- Get principal value
        ZL := POLAR_TO_COMPLEX( L );
        ZR := POLAR_TO_COMPLEX( R );
        ZOUT := COMPLEX_TO_POLAR(COMPLEX'(ZL.RE - ZR.RE, ZL.IM -ZR.IM));
        return ZOUT;
    end "-";

    function "-" ( L: in REAL;  R: in COMPLEX_POLAR) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR'(0.0, 0.0) on error
        --
        variable ZR : COMPLEX;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( R.ARG = -MATH_PI ) then
                assert FALSE
                            report "R.ARG = -MATH_PI in -(L,R)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Get principal value
        ZR := POLAR_TO_COMPLEX( R );
        ZOUT := COMPLEX_TO_POLAR(COMPLEX'(L - ZR.RE, -1.0*ZR.IM));
        return ZOUT;
    end "-";

    function "-" ( L: in COMPLEX_POLAR;  R: in REAL) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR'(0.0, 0.0) on error
        --
        variable ZL : COMPLEX;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( L.ARG = -MATH_PI ) then
                assert FALSE
                            report "L.ARG = -MATH_PI in -(L,R)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Get principal value
        ZL := POLAR_TO_COMPLEX( L );
        ZOUT := COMPLEX_TO_POLAR(COMPLEX'(ZL.RE - R, ZL.IM));
        return ZOUT;
    end "-";


    function "*" ( L: in COMPLEX;  R: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
    begin
        return COMPLEX'(L.RE * R.RE - L.IM * R.IM, L.RE * R.IM + L.IM * R.RE);
    end "*";


    function "*" ( L: in REAL;  R: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
    begin
        return COMPLEX'(L * R.RE, L * R.IM);
    end "*";

    function "*" ( L: in COMPLEX;  R: in REAL )    return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        None
    begin
        return COMPLEX'(L.RE * R, L.IM * R);
    end "*";

    function "*" ( L: in COMPLEX_POLAR; R: in COMPLEX_POLAR)
                                                        return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR'(0.0, 0.0) on error
        --
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( L.ARG = -MATH_PI ) then
                assert FALSE
                            report "L.ARG = -MATH_PI in *(L,R)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        if ( R.ARG = -MATH_PI ) then
                assert FALSE
                            report "R.ARG = -MATH_PI in *(L,R)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Get principal value
        ZOUT.MAG := L.MAG * R.MAG;
        ZOUT.ARG := GET_PRINCIPAL_VALUE(L.ARG + R.ARG);

        return ZOUT;
    end "*";

    function "*" ( L: in REAL;  R: in COMPLEX_POLAR) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR'(0.0, 0.0) on error
        --
            variable ZL : COMPLEX_POLAR;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( R.ARG = -MATH_PI ) then
                assert FALSE
                            report "R.ARG = -MATH_PI in *(L,R)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Get principal value
        ZL.MAG := POSITIVE_REAL'(ABS(L));
        if ( L < 0.0 ) then
                ZL.ARG := MATH_PI;
        else
                ZL.ARG := 0.0;
        end if;

        ZOUT.MAG := ZL.MAG * R.MAG;
        ZOUT.ARG := GET_PRINCIPAL_VALUE(ZL.ARG + R.ARG);

        return ZOUT;
    end "*";

    function "*" ( L: in COMPLEX_POLAR;  R: in REAL) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR'(0.0, 0.0) on error
        --
        variable ZR : COMPLEX_POLAR;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if ( L.ARG = -MATH_PI ) then
                assert FALSE
                            report "L.ARG = -MATH_PI in *(L,R)"
                            severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Get principal value
        ZR.MAG := POSITIVE_REAL'(ABS(R));
        if ( R < 0.0 ) then
                ZR.ARG := MATH_PI;
        else
                ZR.ARG := 0.0;
        end if;

        ZOUT.MAG := L.MAG * ZR.MAG;
        ZOUT.ARG := GET_PRINCIPAL_VALUE(L.ARG + ZR.ARG);

        return ZOUT;
    end "*";

   function "/" ( L: in COMPLEX;  R: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX'(REAL'HIGH, 0.0) on error
        --
        variable TEMP : REAL := R.RE*R.RE + R.IM*R.IM;
   begin
        -- Check validity of input arguments
        if (TEMP = 0.0) then
                 assert FALSE
                        report "Attempt to divide COMPLEX by (0.0, 0.0)"
                        severity ERROR;
                 return COMPLEX'(REAL'HIGH, 0.0);
        end if;

        -- Get value
        return COMPLEX'( (L.RE * R.RE + L.IM * R.IM) / TEMP,
                         (L.IM * R.RE - L.RE * R.IM) / TEMP);
    end "/";

   function "/" ( L: in REAL;  R: in COMPLEX ) return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX'(REAL'HIGH, 0.0) on error
        --
        variable TEMP : REAL := R.RE*R.RE + R.IM*R.IM;
    begin
        -- Check validity of input arguments
        if (TEMP = 0.0) then
                 assert FALSE
                        report "Attempt to divide COMPLEX by (0.0, 0.0)"
                        severity ERROR;
                 return COMPLEX'(REAL'HIGH, 0.0);
        end if;

        -- Get value
        TEMP := L / TEMP;
        return  COMPLEX'( TEMP * R.RE, -TEMP * R.IM );
    end "/";

    function "/" ( L: in COMPLEX;  R: in REAL )    return COMPLEX is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX'(REAL'HIGH, 0.0) on error
    begin
        -- Check validity of input arguments
        if (R = 0.0) then
                 assert FALSE
                        report "Attempt to divide COMPLEX by 0.0"
                        severity ERROR;
                 return COMPLEX'(REAL'HIGH, 0.0);
        end if;

        -- Get value
        return COMPLEX'(L.RE / R, L.IM / R);
    end "/";


    function "/" ( L: in COMPLEX_POLAR; R: in COMPLEX_POLAR)
                                                        return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR'(REAL'HIGH, 0.0) on error
        --
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if (R.MAG = 0.0) then
                assert FALSE
                        report "Attempt to divide COMPLEX_POLAR by (0.0, 0.0)"
                        severity ERROR;
                return COMPLEX_POLAR'(REAL'HIGH, 0.0);
        end if;

        if ( L.ARG = -MATH_PI ) then
                assert FALSE
                        report "L.ARG = -MATH_PI in /(L,R)"
                        severity ERROR;
                return COMPLEX_POLAR'(REAL'HIGH, 0.0);
        end if;

        if ( R.ARG = -MATH_PI ) then
                assert FALSE
                        report "R.ARG = -MATH_PI in /(L,R)"
                        severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Get principal value
        ZOUT.MAG := L.MAG/R.MAG;
        ZOUT.ARG := GET_PRINCIPAL_VALUE(L.ARG - R.ARG);

        return ZOUT;
    end "/";

    function "/" ( L: in COMPLEX_POLAR;  R: in REAL) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR'(REAL'HIGH, 0.0) on error
        --
        variable ZR : COMPLEX_POLAR;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if (R = 0.0) then
                assert FALSE
                        report "Attempt to divide COMPLEX_POLAR by 0.0"
                        severity ERROR;
                return COMPLEX_POLAR'(REAL'HIGH, 0.0);
        end if;

        if ( L.ARG = -MATH_PI ) then
                assert FALSE
                        report "L.ARG = -MATH_PI in /(L,R)"
                        severity ERROR;
                return COMPLEX_POLAR'(REAL'HIGH, 0.0);
        end if;

        -- Get principal value
        ZR.MAG := POSITIVE_REAL'(ABS(R));
        if R < 0.0 then
                ZR.ARG := MATH_PI;
        else
                ZR.ARG := 0.0;
        end if;

        ZOUT.MAG := L.MAG/ZR.MAG;
        ZOUT.ARG := GET_PRINCIPAL_VALUE(L.ARG - ZR.ARG);

        return ZOUT;
    end "/";

    function "/" ( L: in REAL;  R: in COMPLEX_POLAR) return COMPLEX_POLAR is
        -- Description:
        --        See function declaration in IEEE Std 1076.2-1996
        -- Notes:
        --        a) Returns COMPLEX_POLAR'(REAL'HIGH, 0.0) on error
        --
        variable ZL : COMPLEX_POLAR;
        variable ZOUT : COMPLEX_POLAR;
    begin
        -- Check validity of input arguments
        if (R.MAG = 0.0) then
                assert FALSE
                        report "Attempt to divide COMPLEX_POLAR by (0.0, 0.0)"
                        severity ERROR;
                return COMPLEX_POLAR'(REAL'HIGH, 0.0);
        end if;

        if ( R.ARG = -MATH_PI ) then
                assert FALSE
                        report "R.ARG = -MATH_P in /(L,R)"
                        severity ERROR;
                return COMPLEX_POLAR'(0.0, 0.0);
        end if;

        -- Get principal value
        ZL.MAG := POSITIVE_REAL'(ABS(L));
        if L < 0.0 then
                ZL.ARG := MATH_PI;
        else
                ZL.ARG := 0.0;
        end if;

        ZOUT.MAG := ZL.MAG/R.MAG;
        ZOUT.ARG := GET_PRINCIPAL_VALUE(ZL.ARG - R.ARG);

        return ZOUT;
    end "/";

end  MATH_COMPLEX;


-- XSIP watermark, do not delete 67d7842dbbe25473c3c32b93c0da8047785f30d78e8a024de1b57352245f9689
>>>>>>> d68cfb566fed6f983427010d388a4e39e9131875
